/*
 * tt_prim_diode.v
 *
 * TT Primitive
 * Antenna diode
 *
 * Author: Sylvain Munaut <tnt@246tNt.com>
 */

`default_nettype none

module tt_prim_diode (
	inout  wire diode
);

	//pulldown(diode);

endmodule // tt_prim_diode
