magic
tech sky130A
timestamp 1716288850
<< nwell >>
rect 321 2422 470 2558
<< pwell >>
rect 321 2558 470 2684
<< nmos >>
rect 410 2600 425 2642
<< pmoshvt >>
rect 410 2440 425 2540
<< ndiff >>
rect 383 2630 410 2642
rect 383 2612 387 2630
rect 404 2612 410 2630
rect 383 2600 410 2612
rect 425 2630 452 2642
rect 425 2612 431 2630
rect 448 2612 452 2630
rect 425 2600 452 2612
<< pdiff >>
rect 383 2528 410 2540
rect 383 2452 387 2528
rect 404 2452 410 2528
rect 383 2440 410 2452
rect 425 2528 452 2540
rect 425 2452 431 2528
rect 448 2452 452 2528
rect 425 2440 452 2452
<< ndiffc >>
rect 387 2612 404 2630
rect 431 2612 448 2630
<< pdiffc >>
rect 387 2452 404 2528
rect 431 2452 448 2528
<< psubdiff >>
rect 339 2630 356 2642
rect 339 2600 356 2612
<< nsubdiff >>
rect 339 2528 356 2540
rect 339 2440 356 2452
<< psubdiffcont >>
rect 339 2612 356 2630
<< nsubdiffcont >>
rect 339 2452 356 2528
<< poly >>
rect 410 2642 425 2655
rect 410 2586 425 2600
rect 392 2581 425 2586
rect 392 2564 400 2581
rect 417 2564 425 2581
rect 392 2559 425 2564
rect 410 2540 425 2559
rect 410 2427 425 2440
<< polycont >>
rect 400 2564 417 2581
<< locali >>
rect 339 2635 404 2638
rect 339 2630 345 2635
rect 398 2630 404 2635
rect 339 2607 345 2612
rect 398 2607 404 2612
rect 339 2604 404 2607
rect 431 2635 448 2638
rect 431 2604 448 2607
rect 417 2564 425 2581
rect 339 2533 404 2536
rect 339 2528 345 2533
rect 398 2528 404 2533
rect 339 2447 345 2452
rect 398 2447 404 2452
rect 339 2444 404 2447
rect 431 2533 448 2536
rect 431 2444 448 2447
<< viali >>
rect 345 2630 398 2635
rect 345 2612 356 2630
rect 356 2612 387 2630
rect 387 2612 398 2630
rect 345 2607 398 2612
rect 431 2630 448 2635
rect 431 2612 448 2630
rect 431 2607 448 2612
rect 388 2564 400 2581
rect 400 2564 405 2581
rect 345 2528 398 2533
rect 345 2452 356 2528
rect 356 2452 387 2528
rect 387 2452 398 2528
rect 345 2447 398 2452
rect 431 2528 448 2533
rect 431 2452 448 2528
rect 431 2447 448 2452
<< metal1 >>
rect 339 2635 404 2638
rect 339 2607 345 2635
rect 398 2607 404 2635
rect 339 2604 404 2607
rect 425 2635 454 2638
rect 425 2607 431 2635
rect 448 2607 454 2635
rect 382 2581 411 2584
rect 339 2564 388 2581
rect 405 2564 411 2581
rect 382 2561 411 2564
rect 339 2533 404 2536
rect 339 2447 345 2533
rect 398 2447 404 2533
rect 339 2444 404 2447
rect 425 2533 454 2607
rect 425 2447 431 2533
rect 448 2447 454 2533
rect 425 2444 454 2447
<< properties >>
string MASKHINTS_NSDM 326 2550 465 2590
string MASKHINTS_PSDM 326 2550 465 2590
<< end >>
