magic
tech sky130A
magscale 1 2
timestamp 1718533623
<< nwell >>
rect 887 0 2707 670
<< pwell >>
rect 52 0 887 670
<< mvnmos >>
rect 219 363 819 463
rect 219 207 819 307
<< mvpmos >>
rect 953 363 2553 463
rect 953 207 2553 307
<< mvndiff >>
rect 219 508 819 516
rect 219 474 231 508
rect 807 474 819 508
rect 219 463 819 474
rect 219 352 819 363
rect 219 318 231 352
rect 807 318 819 352
rect 219 307 819 318
rect 219 196 819 207
rect 219 162 231 196
rect 807 162 819 196
rect 219 154 819 162
<< mvpdiff >>
rect 953 508 2553 516
rect 953 474 965 508
rect 2541 474 2553 508
rect 953 463 2553 474
rect 953 352 2553 363
rect 953 318 965 352
rect 2541 318 2553 352
rect 953 307 2553 318
rect 953 196 2553 207
rect 953 162 965 196
rect 2541 162 2553 196
rect 953 154 2553 162
<< mvndiffc >>
rect 231 474 807 508
rect 231 318 807 352
rect 231 162 807 196
<< mvpdiffc >>
rect 965 474 2541 508
rect 965 318 2541 352
rect 965 162 2541 196
<< mvpsubdiff >>
rect 111 590 175 624
rect 786 590 810 624
rect 111 560 145 590
rect 111 80 145 110
rect 111 46 175 80
rect 786 46 810 80
<< mvnsubdiff >>
rect 962 570 986 604
rect 2577 570 2641 604
rect 2607 540 2641 570
rect 2607 100 2641 130
rect 962 66 986 100
rect 2577 66 2641 100
<< mvpsubdiffcont >>
rect 175 590 786 624
rect 111 110 145 560
rect 175 46 786 80
<< mvnsubdiffcont >>
rect 986 570 2577 604
rect 2607 130 2641 540
rect 986 66 2577 100
<< poly >>
rect 859 500 913 516
rect 859 463 869 500
rect 193 363 219 463
rect 819 363 869 463
rect 859 307 869 363
rect 193 207 219 307
rect 819 207 869 307
rect 859 170 869 207
rect 903 463 913 500
rect 903 363 953 463
rect 2553 363 2579 463
rect 903 307 913 363
rect 903 207 953 307
rect 2553 207 2579 307
rect 903 170 913 207
rect 859 154 913 170
<< polycont >>
rect 869 170 903 500
<< locali >>
rect 111 590 175 624
rect 795 590 810 624
rect 111 560 145 590
rect 962 570 977 604
rect 2577 570 2641 604
rect 2607 540 2641 570
rect 215 474 231 508
rect 807 474 823 508
rect 869 504 903 516
rect 215 318 231 352
rect 807 318 823 352
rect 215 162 231 196
rect 807 162 823 196
rect 949 474 965 508
rect 2541 474 2557 508
rect 949 318 965 352
rect 2541 318 2557 352
rect 869 154 903 166
rect 949 162 965 196
rect 2541 162 2557 196
rect 111 80 145 110
rect 2607 100 2641 130
rect 111 46 175 80
rect 795 46 810 80
rect 962 66 977 100
rect 2577 66 2641 100
<< viali >>
rect 175 590 786 624
rect 786 590 795 624
rect 977 570 986 604
rect 986 570 2577 604
rect 111 110 145 560
rect 231 474 807 508
rect 869 500 903 504
rect 231 318 807 352
rect 231 162 807 196
rect 869 170 903 500
rect 965 474 2541 508
rect 965 318 2541 352
rect 869 166 903 170
rect 965 162 2541 196
rect 2607 130 2641 540
rect 175 46 786 80
rect 786 46 795 80
rect 977 66 986 100
rect 986 66 2577 100
<< metal1 >>
rect 105 624 819 630
rect 105 590 175 624
rect 795 590 819 624
rect 105 584 819 590
rect 105 560 151 584
rect 105 110 111 560
rect 145 110 151 560
rect 219 508 819 584
rect 953 604 2647 610
rect 953 570 977 604
rect 2577 570 2647 604
rect 953 564 2647 570
rect 219 474 231 508
rect 807 474 819 508
rect 219 468 819 474
rect 860 510 912 516
rect 219 309 225 361
rect 813 309 819 361
rect 105 86 151 110
rect 219 196 819 202
rect 219 162 231 196
rect 807 162 819 196
rect 219 86 819 162
rect 953 508 2553 564
rect 953 474 965 508
rect 2541 474 2553 508
rect 953 468 2553 474
rect 2601 540 2647 564
rect 953 309 959 361
rect 2547 309 2553 361
rect 860 154 912 160
rect 953 196 2553 202
rect 953 162 965 196
rect 2541 162 2553 196
rect 105 80 819 86
rect 105 46 175 80
rect 795 46 819 80
rect 953 106 2553 162
rect 2601 130 2607 540
rect 2641 130 2647 540
rect 2601 106 2647 130
rect 953 100 2647 106
rect 953 66 977 100
rect 2577 66 2647 100
rect 953 60 2647 66
rect 105 40 819 46
<< via1 >>
rect 860 504 912 510
rect 225 352 813 361
rect 225 318 231 352
rect 231 318 807 352
rect 807 318 813 352
rect 225 309 813 318
rect 860 166 869 504
rect 869 166 903 504
rect 903 166 912 504
rect 959 352 2547 361
rect 959 318 965 352
rect 965 318 2541 352
rect 2541 318 2547 352
rect 959 309 2547 318
rect 860 160 912 166
<< metal2 >>
rect 715 568 1057 672
rect 715 361 819 568
rect 219 309 225 361
rect 813 309 819 361
rect 860 510 912 516
rect 953 361 1057 568
rect 953 309 959 361
rect 2547 309 2553 361
rect 860 154 912 160
<< properties >>
string FIXED_BBOX 0 0 2760 670
<< end >>
