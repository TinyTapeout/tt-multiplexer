magic
tech sky130A
magscale 1 2
timestamp 1718439036
<< nwell >>
rect 594 0 1827 644
<< pwell >>
rect 13 0 594 644
<< nmos >>
rect 160 437 510 467
rect 160 351 510 381
rect 160 263 510 293
rect 160 177 510 207
<< pmoshvt >>
rect 630 437 1680 467
rect 630 351 1680 381
rect 630 263 1680 293
rect 630 177 1680 207
<< ndiff >>
rect 160 512 510 520
rect 160 478 172 512
rect 498 478 510 512
rect 160 467 510 478
rect 160 426 510 437
rect 160 392 172 426
rect 498 392 510 426
rect 160 381 510 392
rect 160 338 510 351
rect 160 304 172 338
rect 498 304 510 338
rect 160 293 510 304
rect 160 252 510 263
rect 160 218 172 252
rect 498 218 510 252
rect 160 207 510 218
rect 160 166 510 177
rect 160 132 172 166
rect 498 132 510 166
rect 160 124 510 132
<< pdiff >>
rect 630 512 1680 520
rect 630 478 642 512
rect 1668 478 1680 512
rect 630 467 1680 478
rect 630 426 1680 437
rect 630 392 642 426
rect 1668 392 1680 426
rect 630 381 1680 392
rect 630 338 1680 351
rect 630 304 642 338
rect 1668 304 1680 338
rect 630 293 1680 304
rect 630 252 1680 263
rect 630 218 642 252
rect 1668 218 1680 252
rect 630 207 1680 218
rect 630 166 1680 177
rect 630 132 642 166
rect 1668 132 1680 166
rect 630 124 1680 132
<< ndiffc >>
rect 172 478 498 512
rect 172 392 498 426
rect 172 304 498 338
rect 172 218 498 252
rect 172 132 498 166
<< pdiffc >>
rect 642 478 1668 512
rect 642 392 1668 426
rect 642 304 1668 338
rect 642 218 1668 252
rect 642 132 1668 166
<< psubdiff >>
rect 72 574 136 608
rect 480 574 504 608
rect 72 544 106 574
rect 72 70 106 100
rect 72 36 136 70
rect 480 36 504 70
<< nsubdiff >>
rect 636 574 660 608
rect 1704 574 1768 608
rect 1734 544 1768 574
rect 1734 70 1768 100
rect 636 36 660 70
rect 1704 36 1768 70
<< psubdiffcont >>
rect 136 574 480 608
rect 72 100 106 544
rect 136 36 480 70
<< nsubdiffcont >>
rect 660 574 1704 608
rect 1734 100 1768 544
rect 660 36 1704 70
<< poly >>
rect 538 504 592 520
rect 538 467 548 504
rect 134 437 160 467
rect 510 437 548 467
rect 538 381 548 437
rect 134 351 160 381
rect 510 351 548 381
rect 538 293 548 351
rect 134 263 160 293
rect 510 263 548 293
rect 538 207 548 263
rect 134 177 160 207
rect 510 177 548 207
rect 538 140 548 177
rect 582 467 592 504
rect 582 437 630 467
rect 1680 437 1706 467
rect 582 381 592 437
rect 582 351 630 381
rect 1680 351 1706 381
rect 582 293 592 351
rect 582 263 630 293
rect 1680 263 1706 293
rect 582 207 592 263
rect 582 177 630 207
rect 1680 177 1706 207
rect 582 140 592 177
rect 538 124 592 140
<< polycont >>
rect 548 140 582 504
<< locali >>
rect 72 574 136 608
rect 480 574 510 608
rect 630 574 660 608
rect 1704 574 1768 608
rect 72 544 106 574
rect 1734 544 1768 574
rect 156 478 172 512
rect 498 478 514 512
rect 548 504 550 520
rect 156 392 172 426
rect 498 392 514 426
rect 156 304 172 338
rect 498 304 514 338
rect 156 218 172 252
rect 498 218 514 252
rect 156 132 172 166
rect 498 132 514 166
rect 548 124 550 140
rect 590 124 592 520
rect 626 478 642 512
rect 1668 478 1684 512
rect 626 392 642 426
rect 1668 392 1684 426
rect 626 304 642 338
rect 1668 304 1684 338
rect 626 218 642 252
rect 1668 218 1684 252
rect 626 132 642 166
rect 1668 132 1684 166
rect 72 70 106 100
rect 1734 70 1768 100
rect 72 36 136 70
rect 480 36 510 70
rect 630 36 660 70
rect 1704 36 1768 70
<< viali >>
rect 136 574 480 608
rect 660 574 1704 608
rect 72 100 106 544
rect 172 478 498 512
rect 550 504 590 520
rect 172 392 498 426
rect 172 304 498 338
rect 172 218 498 252
rect 172 132 498 166
rect 550 140 582 504
rect 582 140 590 504
rect 550 124 590 140
rect 642 478 1668 512
rect 642 392 1668 426
rect 642 304 1668 338
rect 642 218 1668 252
rect 642 132 1668 166
rect 1734 100 1768 544
rect 136 36 480 70
rect 660 36 1704 70
<< metal1 >>
rect 66 608 166 614
rect 366 608 510 614
rect 66 574 136 608
rect 480 574 510 608
rect 66 568 166 574
rect 66 544 112 568
rect 66 100 72 544
rect 106 348 112 544
rect 160 472 166 568
rect 366 512 510 574
rect 630 608 774 614
rect 1674 608 1774 614
rect 630 574 660 608
rect 1704 574 1774 608
rect 498 478 510 512
rect 366 472 510 478
rect 544 526 596 532
rect 160 383 166 435
rect 504 383 510 435
rect 366 346 372 348
rect 366 338 510 346
rect 498 304 510 338
rect 366 298 510 304
rect 366 296 372 298
rect 106 100 112 296
rect 160 209 166 261
rect 504 209 510 261
rect 66 76 112 100
rect 160 76 166 172
rect 66 70 166 76
rect 66 36 136 70
rect 66 30 166 36
rect 504 30 510 172
rect 630 512 774 574
rect 1674 568 1774 574
rect 630 478 642 512
rect 630 472 774 478
rect 1674 472 1680 568
rect 1728 544 1774 568
rect 630 383 636 435
rect 1674 383 1680 435
rect 1728 348 1734 544
rect 768 346 774 348
rect 630 338 774 346
rect 630 304 642 338
rect 630 298 774 304
rect 768 296 774 298
rect 630 209 636 261
rect 1674 209 1680 261
rect 544 112 596 118
rect 630 30 636 172
rect 1674 76 1680 172
rect 1728 100 1734 296
rect 1768 100 1774 544
rect 1728 76 1774 100
rect 1674 70 1774 76
rect 1704 36 1774 70
rect 1674 30 1774 36
<< via1 >>
rect 166 608 366 614
rect 166 574 366 608
rect 166 512 366 574
rect 774 608 1674 614
rect 774 574 1674 608
rect 166 478 172 512
rect 172 478 366 512
rect 166 472 366 478
rect 544 520 596 526
rect 166 426 504 435
rect 166 392 172 426
rect 172 392 498 426
rect 498 392 504 426
rect 166 383 504 392
rect 72 296 106 348
rect 106 338 366 348
rect 106 304 172 338
rect 172 304 366 338
rect 106 296 366 304
rect 166 252 504 261
rect 166 218 172 252
rect 172 218 498 252
rect 498 218 504 252
rect 166 209 504 218
rect 166 166 504 172
rect 166 132 172 166
rect 172 132 498 166
rect 498 132 504 166
rect 166 70 504 132
rect 166 36 480 70
rect 480 36 504 70
rect 166 30 504 36
rect 544 124 550 520
rect 550 124 590 520
rect 590 124 596 520
rect 774 512 1674 574
rect 774 478 1668 512
rect 1668 478 1674 512
rect 774 472 1674 478
rect 636 426 1674 435
rect 636 392 642 426
rect 642 392 1668 426
rect 1668 392 1674 426
rect 636 383 1674 392
rect 774 338 1734 348
rect 774 304 1668 338
rect 1668 304 1734 338
rect 774 296 1734 304
rect 1734 296 1768 348
rect 636 252 1674 261
rect 636 218 642 252
rect 642 218 1668 252
rect 1668 218 1674 252
rect 636 209 1674 218
rect 544 118 596 124
rect 636 166 1674 172
rect 636 132 642 166
rect 642 132 1668 166
rect 1668 132 1674 166
rect 636 70 1674 132
rect 636 36 660 70
rect 660 36 1674 70
rect 636 30 1674 36
<< metal2 >>
rect 66 472 166 614
rect 366 472 372 614
rect 406 566 734 644
rect 66 348 126 472
rect 406 435 510 566
rect 160 383 166 435
rect 504 383 510 435
rect 66 296 72 348
rect 366 296 372 348
rect 66 172 126 296
rect 406 261 510 383
rect 160 209 166 261
rect 504 209 510 261
rect 544 526 596 532
rect 66 30 166 172
rect 504 30 510 172
rect 630 435 734 566
rect 768 472 774 614
rect 1674 472 1774 614
rect 630 383 636 435
rect 1674 383 1680 435
rect 630 261 734 383
rect 1714 348 1774 472
rect 768 296 774 348
rect 1768 296 1774 348
rect 630 209 636 261
rect 1674 209 1680 261
rect 1714 172 1774 296
rect 544 0 596 118
rect 630 30 636 172
rect 1674 30 1774 172
<< properties >>
string FIXED_BBOX 0 0 1840 644
<< end >>
