magic
tech sky130A
magscale 1 2
timestamp 1520178628
<< checkpaint >>
rect -1239 -1240 10328 16120
<< metal3 >>
rect 21 14832 9060 14860
rect 21 10128 29 14832
rect 4013 10128 9060 14832
rect 21 10060 9060 10128
rect 4501 9742 9063 9770
rect 4501 5198 4509 9742
rect 8493 5198 9063 9742
rect 4501 5108 9063 5198
rect 21 4787 9068 4809
rect 21 83 29 4787
rect 4013 83 9068 4787
rect 21 20 9068 83
<< via3 >>
rect 29 10128 4013 14832
rect 4509 5198 8493 9742
rect 29 83 4013 4787
<< properties >>
string FIXED_BBOX 0 0 9080 14920
<< end >>
