magic
tech sky130A
magscale 1 2
timestamp 1709841855
<< nwell >>
rect 0 490 1838 21944
<< pmos >>
rect 219 21714 1619 21744
rect 219 21618 1619 21648
rect 219 21522 1619 21552
rect 219 21426 1619 21456
rect 219 21330 1619 21360
rect 219 21234 1619 21264
rect 219 21138 1619 21168
rect 219 21042 1619 21072
rect 219 20946 1619 20976
rect 219 20850 1619 20880
rect 219 20754 1619 20784
rect 219 20658 1619 20688
rect 219 20562 1619 20592
rect 219 20466 1619 20496
rect 219 20370 1619 20400
rect 219 20274 1619 20304
rect 219 20178 1619 20208
rect 219 20082 1619 20112
rect 219 19986 1619 20016
rect 219 19890 1619 19920
rect 219 19794 1619 19824
rect 219 19698 1619 19728
rect 219 19602 1619 19632
rect 219 19506 1619 19536
rect 219 19410 1619 19440
rect 219 19314 1619 19344
rect 219 19218 1619 19248
rect 219 19122 1619 19152
rect 219 19026 1619 19056
rect 219 18930 1619 18960
rect 219 18834 1619 18864
rect 219 18738 1619 18768
rect 219 18642 1619 18672
rect 219 18546 1619 18576
rect 219 18450 1619 18480
rect 219 18354 1619 18384
rect 219 18258 1619 18288
rect 219 18162 1619 18192
rect 219 18066 1619 18096
rect 219 17970 1619 18000
rect 219 17874 1619 17904
rect 219 17778 1619 17808
rect 219 17682 1619 17712
rect 219 17586 1619 17616
rect 219 17490 1619 17520
rect 219 17394 1619 17424
rect 219 17298 1619 17328
rect 219 17202 1619 17232
rect 219 17106 1619 17136
rect 219 17010 1619 17040
rect 219 16914 1619 16944
rect 219 16818 1619 16848
rect 219 16722 1619 16752
rect 219 16626 1619 16656
rect 219 16530 1619 16560
rect 219 16434 1619 16464
rect 219 16338 1619 16368
rect 219 16242 1619 16272
rect 219 16146 1619 16176
rect 219 16050 1619 16080
rect 219 15954 1619 15984
rect 219 15858 1619 15888
rect 219 15762 1619 15792
rect 219 15666 1619 15696
rect 219 15570 1619 15600
rect 219 15474 1619 15504
rect 219 15378 1619 15408
rect 219 15282 1619 15312
rect 219 15186 1619 15216
rect 219 15090 1619 15120
rect 219 14994 1619 15024
rect 219 14898 1619 14928
rect 219 14802 1619 14832
rect 219 14706 1619 14736
rect 219 14610 1619 14640
rect 219 14514 1619 14544
rect 219 14418 1619 14448
rect 219 14322 1619 14352
rect 219 14226 1619 14256
rect 219 14130 1619 14160
rect 219 14034 1619 14064
rect 219 13938 1619 13968
rect 219 13842 1619 13872
rect 219 13746 1619 13776
rect 219 13650 1619 13680
rect 219 13554 1619 13584
rect 219 13458 1619 13488
rect 219 13362 1619 13392
rect 219 13266 1619 13296
rect 219 13170 1619 13200
rect 219 13074 1619 13104
rect 219 12978 1619 13008
rect 219 12882 1619 12912
rect 219 12786 1619 12816
rect 219 12690 1619 12720
rect 219 12594 1619 12624
rect 219 12498 1619 12528
rect 219 12402 1619 12432
rect 219 12306 1619 12336
rect 219 12210 1619 12240
rect 219 12114 1619 12144
rect 219 12018 1619 12048
rect 219 11922 1619 11952
rect 219 11826 1619 11856
rect 219 11730 1619 11760
rect 219 11634 1619 11664
rect 219 11538 1619 11568
rect 219 11442 1619 11472
rect 219 11346 1619 11376
rect 219 11250 1619 11280
rect 219 11154 1619 11184
rect 219 11058 1619 11088
rect 219 10962 1619 10992
rect 219 10866 1619 10896
rect 219 10770 1619 10800
rect 219 10674 1619 10704
rect 219 10578 1619 10608
rect 219 10482 1619 10512
rect 219 10386 1619 10416
rect 219 10290 1619 10320
rect 219 10194 1619 10224
rect 219 10098 1619 10128
rect 219 10002 1619 10032
rect 219 9906 1619 9936
rect 219 9810 1619 9840
rect 219 9714 1619 9744
rect 219 9618 1619 9648
rect 219 9522 1619 9552
rect 219 9426 1619 9456
rect 219 9330 1619 9360
rect 219 9234 1619 9264
rect 219 9138 1619 9168
rect 219 9042 1619 9072
rect 219 8946 1619 8976
rect 219 8850 1619 8880
rect 219 8754 1619 8784
rect 219 8658 1619 8688
rect 219 8562 1619 8592
rect 219 8466 1619 8496
rect 219 8370 1619 8400
rect 219 8274 1619 8304
rect 219 8178 1619 8208
rect 219 8082 1619 8112
rect 219 7986 1619 8016
rect 219 7890 1619 7920
rect 219 7794 1619 7824
rect 219 7698 1619 7728
rect 219 7602 1619 7632
rect 219 7506 1619 7536
rect 219 7410 1619 7440
rect 219 7314 1619 7344
rect 219 7218 1619 7248
rect 219 7122 1619 7152
rect 219 7026 1619 7056
rect 219 6930 1619 6960
rect 219 6834 1619 6864
rect 219 6738 1619 6768
rect 219 6642 1619 6672
rect 219 6546 1619 6576
rect 219 6450 1619 6480
rect 219 6354 1619 6384
rect 219 6258 1619 6288
rect 219 6162 1619 6192
rect 219 6066 1619 6096
rect 219 5970 1619 6000
rect 219 5874 1619 5904
rect 219 5778 1619 5808
rect 219 5682 1619 5712
rect 219 5586 1619 5616
rect 219 5490 1619 5520
rect 219 5394 1619 5424
rect 219 5298 1619 5328
rect 219 5202 1619 5232
rect 219 5106 1619 5136
rect 219 5010 1619 5040
rect 219 4914 1619 4944
rect 219 4818 1619 4848
rect 219 4722 1619 4752
rect 219 4626 1619 4656
rect 219 4530 1619 4560
rect 219 4434 1619 4464
rect 219 4338 1619 4368
rect 219 4242 1619 4272
rect 219 4146 1619 4176
rect 219 4050 1619 4080
rect 219 3954 1619 3984
rect 219 3858 1619 3888
rect 219 3762 1619 3792
rect 219 3666 1619 3696
rect 219 3570 1619 3600
rect 219 3474 1619 3504
rect 219 3378 1619 3408
rect 219 3282 1619 3312
rect 219 3186 1619 3216
rect 219 3090 1619 3120
rect 219 2994 1619 3024
rect 219 2898 1619 2928
rect 219 2802 1619 2832
rect 219 2706 1619 2736
rect 219 2610 1619 2640
rect 219 2514 1619 2544
rect 219 2418 1619 2448
rect 219 2322 1619 2352
rect 219 2226 1619 2256
rect 219 2130 1619 2160
rect 219 2034 1619 2064
rect 219 1938 1619 1968
rect 219 1842 1619 1872
rect 219 1746 1619 1776
rect 219 1650 1619 1680
rect 219 1554 1619 1584
rect 219 1458 1619 1488
rect 219 1362 1619 1392
rect 219 1266 1619 1296
rect 219 1170 1619 1200
rect 219 1074 1619 1104
rect 219 978 1619 1008
rect 219 882 1619 912
rect 219 786 1619 816
rect 219 690 1619 720
<< pdiff >>
rect 219 21794 1619 21806
rect 219 21760 231 21794
rect 1607 21760 1619 21794
rect 219 21744 1619 21760
rect 219 21698 1619 21714
rect 219 21664 231 21698
rect 1607 21664 1619 21698
rect 219 21648 1619 21664
rect 219 21602 1619 21618
rect 219 21568 231 21602
rect 1607 21568 1619 21602
rect 219 21552 1619 21568
rect 219 21506 1619 21522
rect 219 21472 231 21506
rect 1607 21472 1619 21506
rect 219 21456 1619 21472
rect 219 21410 1619 21426
rect 219 21376 231 21410
rect 1607 21376 1619 21410
rect 219 21360 1619 21376
rect 219 21314 1619 21330
rect 219 21280 231 21314
rect 1607 21280 1619 21314
rect 219 21264 1619 21280
rect 219 21218 1619 21234
rect 219 21184 231 21218
rect 1607 21184 1619 21218
rect 219 21168 1619 21184
rect 219 21122 1619 21138
rect 219 21088 231 21122
rect 1607 21088 1619 21122
rect 219 21072 1619 21088
rect 219 21026 1619 21042
rect 219 20992 231 21026
rect 1607 20992 1619 21026
rect 219 20976 1619 20992
rect 219 20930 1619 20946
rect 219 20896 231 20930
rect 1607 20896 1619 20930
rect 219 20880 1619 20896
rect 219 20834 1619 20850
rect 219 20800 231 20834
rect 1607 20800 1619 20834
rect 219 20784 1619 20800
rect 219 20738 1619 20754
rect 219 20704 231 20738
rect 1607 20704 1619 20738
rect 219 20688 1619 20704
rect 219 20642 1619 20658
rect 219 20608 231 20642
rect 1607 20608 1619 20642
rect 219 20592 1619 20608
rect 219 20546 1619 20562
rect 219 20512 231 20546
rect 1607 20512 1619 20546
rect 219 20496 1619 20512
rect 219 20450 1619 20466
rect 219 20416 231 20450
rect 1607 20416 1619 20450
rect 219 20400 1619 20416
rect 219 20354 1619 20370
rect 219 20320 231 20354
rect 1607 20320 1619 20354
rect 219 20304 1619 20320
rect 219 20258 1619 20274
rect 219 20224 231 20258
rect 1607 20224 1619 20258
rect 219 20208 1619 20224
rect 219 20162 1619 20178
rect 219 20128 231 20162
rect 1607 20128 1619 20162
rect 219 20112 1619 20128
rect 219 20066 1619 20082
rect 219 20032 231 20066
rect 1607 20032 1619 20066
rect 219 20016 1619 20032
rect 219 19970 1619 19986
rect 219 19936 231 19970
rect 1607 19936 1619 19970
rect 219 19920 1619 19936
rect 219 19874 1619 19890
rect 219 19840 231 19874
rect 1607 19840 1619 19874
rect 219 19824 1619 19840
rect 219 19778 1619 19794
rect 219 19744 231 19778
rect 1607 19744 1619 19778
rect 219 19728 1619 19744
rect 219 19682 1619 19698
rect 219 19648 231 19682
rect 1607 19648 1619 19682
rect 219 19632 1619 19648
rect 219 19586 1619 19602
rect 219 19552 231 19586
rect 1607 19552 1619 19586
rect 219 19536 1619 19552
rect 219 19490 1619 19506
rect 219 19456 231 19490
rect 1607 19456 1619 19490
rect 219 19440 1619 19456
rect 219 19394 1619 19410
rect 219 19360 231 19394
rect 1607 19360 1619 19394
rect 219 19344 1619 19360
rect 219 19298 1619 19314
rect 219 19264 231 19298
rect 1607 19264 1619 19298
rect 219 19248 1619 19264
rect 219 19202 1619 19218
rect 219 19168 231 19202
rect 1607 19168 1619 19202
rect 219 19152 1619 19168
rect 219 19106 1619 19122
rect 219 19072 231 19106
rect 1607 19072 1619 19106
rect 219 19056 1619 19072
rect 219 19010 1619 19026
rect 219 18976 231 19010
rect 1607 18976 1619 19010
rect 219 18960 1619 18976
rect 219 18914 1619 18930
rect 219 18880 231 18914
rect 1607 18880 1619 18914
rect 219 18864 1619 18880
rect 219 18818 1619 18834
rect 219 18784 231 18818
rect 1607 18784 1619 18818
rect 219 18768 1619 18784
rect 219 18722 1619 18738
rect 219 18688 231 18722
rect 1607 18688 1619 18722
rect 219 18672 1619 18688
rect 219 18626 1619 18642
rect 219 18592 231 18626
rect 1607 18592 1619 18626
rect 219 18576 1619 18592
rect 219 18530 1619 18546
rect 219 18496 231 18530
rect 1607 18496 1619 18530
rect 219 18480 1619 18496
rect 219 18434 1619 18450
rect 219 18400 231 18434
rect 1607 18400 1619 18434
rect 219 18384 1619 18400
rect 219 18338 1619 18354
rect 219 18304 231 18338
rect 1607 18304 1619 18338
rect 219 18288 1619 18304
rect 219 18242 1619 18258
rect 219 18208 231 18242
rect 1607 18208 1619 18242
rect 219 18192 1619 18208
rect 219 18146 1619 18162
rect 219 18112 231 18146
rect 1607 18112 1619 18146
rect 219 18096 1619 18112
rect 219 18050 1619 18066
rect 219 18016 231 18050
rect 1607 18016 1619 18050
rect 219 18000 1619 18016
rect 219 17954 1619 17970
rect 219 17920 231 17954
rect 1607 17920 1619 17954
rect 219 17904 1619 17920
rect 219 17858 1619 17874
rect 219 17824 231 17858
rect 1607 17824 1619 17858
rect 219 17808 1619 17824
rect 219 17762 1619 17778
rect 219 17728 231 17762
rect 1607 17728 1619 17762
rect 219 17712 1619 17728
rect 219 17666 1619 17682
rect 219 17632 231 17666
rect 1607 17632 1619 17666
rect 219 17616 1619 17632
rect 219 17570 1619 17586
rect 219 17536 231 17570
rect 1607 17536 1619 17570
rect 219 17520 1619 17536
rect 219 17474 1619 17490
rect 219 17440 231 17474
rect 1607 17440 1619 17474
rect 219 17424 1619 17440
rect 219 17378 1619 17394
rect 219 17344 231 17378
rect 1607 17344 1619 17378
rect 219 17328 1619 17344
rect 219 17282 1619 17298
rect 219 17248 231 17282
rect 1607 17248 1619 17282
rect 219 17232 1619 17248
rect 219 17186 1619 17202
rect 219 17152 231 17186
rect 1607 17152 1619 17186
rect 219 17136 1619 17152
rect 219 17090 1619 17106
rect 219 17056 231 17090
rect 1607 17056 1619 17090
rect 219 17040 1619 17056
rect 219 16994 1619 17010
rect 219 16960 231 16994
rect 1607 16960 1619 16994
rect 219 16944 1619 16960
rect 219 16898 1619 16914
rect 219 16864 231 16898
rect 1607 16864 1619 16898
rect 219 16848 1619 16864
rect 219 16802 1619 16818
rect 219 16768 231 16802
rect 1607 16768 1619 16802
rect 219 16752 1619 16768
rect 219 16706 1619 16722
rect 219 16672 231 16706
rect 1607 16672 1619 16706
rect 219 16656 1619 16672
rect 219 16610 1619 16626
rect 219 16576 231 16610
rect 1607 16576 1619 16610
rect 219 16560 1619 16576
rect 219 16514 1619 16530
rect 219 16480 231 16514
rect 1607 16480 1619 16514
rect 219 16464 1619 16480
rect 219 16418 1619 16434
rect 219 16384 231 16418
rect 1607 16384 1619 16418
rect 219 16368 1619 16384
rect 219 16322 1619 16338
rect 219 16288 231 16322
rect 1607 16288 1619 16322
rect 219 16272 1619 16288
rect 219 16226 1619 16242
rect 219 16192 231 16226
rect 1607 16192 1619 16226
rect 219 16176 1619 16192
rect 219 16130 1619 16146
rect 219 16096 231 16130
rect 1607 16096 1619 16130
rect 219 16080 1619 16096
rect 219 16034 1619 16050
rect 219 16000 231 16034
rect 1607 16000 1619 16034
rect 219 15984 1619 16000
rect 219 15938 1619 15954
rect 219 15904 231 15938
rect 1607 15904 1619 15938
rect 219 15888 1619 15904
rect 219 15842 1619 15858
rect 219 15808 231 15842
rect 1607 15808 1619 15842
rect 219 15792 1619 15808
rect 219 15746 1619 15762
rect 219 15712 231 15746
rect 1607 15712 1619 15746
rect 219 15696 1619 15712
rect 219 15650 1619 15666
rect 219 15616 231 15650
rect 1607 15616 1619 15650
rect 219 15600 1619 15616
rect 219 15554 1619 15570
rect 219 15520 231 15554
rect 1607 15520 1619 15554
rect 219 15504 1619 15520
rect 219 15458 1619 15474
rect 219 15424 231 15458
rect 1607 15424 1619 15458
rect 219 15408 1619 15424
rect 219 15362 1619 15378
rect 219 15328 231 15362
rect 1607 15328 1619 15362
rect 219 15312 1619 15328
rect 219 15266 1619 15282
rect 219 15232 231 15266
rect 1607 15232 1619 15266
rect 219 15216 1619 15232
rect 219 15170 1619 15186
rect 219 15136 231 15170
rect 1607 15136 1619 15170
rect 219 15120 1619 15136
rect 219 15074 1619 15090
rect 219 15040 231 15074
rect 1607 15040 1619 15074
rect 219 15024 1619 15040
rect 219 14978 1619 14994
rect 219 14944 231 14978
rect 1607 14944 1619 14978
rect 219 14928 1619 14944
rect 219 14882 1619 14898
rect 219 14848 231 14882
rect 1607 14848 1619 14882
rect 219 14832 1619 14848
rect 219 14786 1619 14802
rect 219 14752 231 14786
rect 1607 14752 1619 14786
rect 219 14736 1619 14752
rect 219 14690 1619 14706
rect 219 14656 231 14690
rect 1607 14656 1619 14690
rect 219 14640 1619 14656
rect 219 14594 1619 14610
rect 219 14560 231 14594
rect 1607 14560 1619 14594
rect 219 14544 1619 14560
rect 219 14498 1619 14514
rect 219 14464 231 14498
rect 1607 14464 1619 14498
rect 219 14448 1619 14464
rect 219 14402 1619 14418
rect 219 14368 231 14402
rect 1607 14368 1619 14402
rect 219 14352 1619 14368
rect 219 14306 1619 14322
rect 219 14272 231 14306
rect 1607 14272 1619 14306
rect 219 14256 1619 14272
rect 219 14210 1619 14226
rect 219 14176 231 14210
rect 1607 14176 1619 14210
rect 219 14160 1619 14176
rect 219 14114 1619 14130
rect 219 14080 231 14114
rect 1607 14080 1619 14114
rect 219 14064 1619 14080
rect 219 14018 1619 14034
rect 219 13984 231 14018
rect 1607 13984 1619 14018
rect 219 13968 1619 13984
rect 219 13922 1619 13938
rect 219 13888 231 13922
rect 1607 13888 1619 13922
rect 219 13872 1619 13888
rect 219 13826 1619 13842
rect 219 13792 231 13826
rect 1607 13792 1619 13826
rect 219 13776 1619 13792
rect 219 13730 1619 13746
rect 219 13696 231 13730
rect 1607 13696 1619 13730
rect 219 13680 1619 13696
rect 219 13634 1619 13650
rect 219 13600 231 13634
rect 1607 13600 1619 13634
rect 219 13584 1619 13600
rect 219 13538 1619 13554
rect 219 13504 231 13538
rect 1607 13504 1619 13538
rect 219 13488 1619 13504
rect 219 13442 1619 13458
rect 219 13408 231 13442
rect 1607 13408 1619 13442
rect 219 13392 1619 13408
rect 219 13346 1619 13362
rect 219 13312 231 13346
rect 1607 13312 1619 13346
rect 219 13296 1619 13312
rect 219 13250 1619 13266
rect 219 13216 231 13250
rect 1607 13216 1619 13250
rect 219 13200 1619 13216
rect 219 13154 1619 13170
rect 219 13120 231 13154
rect 1607 13120 1619 13154
rect 219 13104 1619 13120
rect 219 13058 1619 13074
rect 219 13024 231 13058
rect 1607 13024 1619 13058
rect 219 13008 1619 13024
rect 219 12962 1619 12978
rect 219 12928 231 12962
rect 1607 12928 1619 12962
rect 219 12912 1619 12928
rect 219 12866 1619 12882
rect 219 12832 231 12866
rect 1607 12832 1619 12866
rect 219 12816 1619 12832
rect 219 12770 1619 12786
rect 219 12736 231 12770
rect 1607 12736 1619 12770
rect 219 12720 1619 12736
rect 219 12674 1619 12690
rect 219 12640 231 12674
rect 1607 12640 1619 12674
rect 219 12624 1619 12640
rect 219 12578 1619 12594
rect 219 12544 231 12578
rect 1607 12544 1619 12578
rect 219 12528 1619 12544
rect 219 12482 1619 12498
rect 219 12448 231 12482
rect 1607 12448 1619 12482
rect 219 12432 1619 12448
rect 219 12386 1619 12402
rect 219 12352 231 12386
rect 1607 12352 1619 12386
rect 219 12336 1619 12352
rect 219 12290 1619 12306
rect 219 12256 231 12290
rect 1607 12256 1619 12290
rect 219 12240 1619 12256
rect 219 12194 1619 12210
rect 219 12160 231 12194
rect 1607 12160 1619 12194
rect 219 12144 1619 12160
rect 219 12098 1619 12114
rect 219 12064 231 12098
rect 1607 12064 1619 12098
rect 219 12048 1619 12064
rect 219 12002 1619 12018
rect 219 11968 231 12002
rect 1607 11968 1619 12002
rect 219 11952 1619 11968
rect 219 11906 1619 11922
rect 219 11872 231 11906
rect 1607 11872 1619 11906
rect 219 11856 1619 11872
rect 219 11810 1619 11826
rect 219 11776 231 11810
rect 1607 11776 1619 11810
rect 219 11760 1619 11776
rect 219 11714 1619 11730
rect 219 11680 231 11714
rect 1607 11680 1619 11714
rect 219 11664 1619 11680
rect 219 11618 1619 11634
rect 219 11584 231 11618
rect 1607 11584 1619 11618
rect 219 11568 1619 11584
rect 219 11522 1619 11538
rect 219 11488 231 11522
rect 1607 11488 1619 11522
rect 219 11472 1619 11488
rect 219 11426 1619 11442
rect 219 11392 231 11426
rect 1607 11392 1619 11426
rect 219 11376 1619 11392
rect 219 11330 1619 11346
rect 219 11296 231 11330
rect 1607 11296 1619 11330
rect 219 11280 1619 11296
rect 219 11234 1619 11250
rect 219 11200 231 11234
rect 1607 11200 1619 11234
rect 219 11184 1619 11200
rect 219 11138 1619 11154
rect 219 11104 231 11138
rect 1607 11104 1619 11138
rect 219 11088 1619 11104
rect 219 11042 1619 11058
rect 219 11008 231 11042
rect 1607 11008 1619 11042
rect 219 10992 1619 11008
rect 219 10946 1619 10962
rect 219 10912 231 10946
rect 1607 10912 1619 10946
rect 219 10896 1619 10912
rect 219 10850 1619 10866
rect 219 10816 231 10850
rect 1607 10816 1619 10850
rect 219 10800 1619 10816
rect 219 10754 1619 10770
rect 219 10720 231 10754
rect 1607 10720 1619 10754
rect 219 10704 1619 10720
rect 219 10658 1619 10674
rect 219 10624 231 10658
rect 1607 10624 1619 10658
rect 219 10608 1619 10624
rect 219 10562 1619 10578
rect 219 10528 231 10562
rect 1607 10528 1619 10562
rect 219 10512 1619 10528
rect 219 10466 1619 10482
rect 219 10432 231 10466
rect 1607 10432 1619 10466
rect 219 10416 1619 10432
rect 219 10370 1619 10386
rect 219 10336 231 10370
rect 1607 10336 1619 10370
rect 219 10320 1619 10336
rect 219 10274 1619 10290
rect 219 10240 231 10274
rect 1607 10240 1619 10274
rect 219 10224 1619 10240
rect 219 10178 1619 10194
rect 219 10144 231 10178
rect 1607 10144 1619 10178
rect 219 10128 1619 10144
rect 219 10082 1619 10098
rect 219 10048 231 10082
rect 1607 10048 1619 10082
rect 219 10032 1619 10048
rect 219 9986 1619 10002
rect 219 9952 231 9986
rect 1607 9952 1619 9986
rect 219 9936 1619 9952
rect 219 9890 1619 9906
rect 219 9856 231 9890
rect 1607 9856 1619 9890
rect 219 9840 1619 9856
rect 219 9794 1619 9810
rect 219 9760 231 9794
rect 1607 9760 1619 9794
rect 219 9744 1619 9760
rect 219 9698 1619 9714
rect 219 9664 231 9698
rect 1607 9664 1619 9698
rect 219 9648 1619 9664
rect 219 9602 1619 9618
rect 219 9568 231 9602
rect 1607 9568 1619 9602
rect 219 9552 1619 9568
rect 219 9506 1619 9522
rect 219 9472 231 9506
rect 1607 9472 1619 9506
rect 219 9456 1619 9472
rect 219 9410 1619 9426
rect 219 9376 231 9410
rect 1607 9376 1619 9410
rect 219 9360 1619 9376
rect 219 9314 1619 9330
rect 219 9280 231 9314
rect 1607 9280 1619 9314
rect 219 9264 1619 9280
rect 219 9218 1619 9234
rect 219 9184 231 9218
rect 1607 9184 1619 9218
rect 219 9168 1619 9184
rect 219 9122 1619 9138
rect 219 9088 231 9122
rect 1607 9088 1619 9122
rect 219 9072 1619 9088
rect 219 9026 1619 9042
rect 219 8992 231 9026
rect 1607 8992 1619 9026
rect 219 8976 1619 8992
rect 219 8930 1619 8946
rect 219 8896 231 8930
rect 1607 8896 1619 8930
rect 219 8880 1619 8896
rect 219 8834 1619 8850
rect 219 8800 231 8834
rect 1607 8800 1619 8834
rect 219 8784 1619 8800
rect 219 8738 1619 8754
rect 219 8704 231 8738
rect 1607 8704 1619 8738
rect 219 8688 1619 8704
rect 219 8642 1619 8658
rect 219 8608 231 8642
rect 1607 8608 1619 8642
rect 219 8592 1619 8608
rect 219 8546 1619 8562
rect 219 8512 231 8546
rect 1607 8512 1619 8546
rect 219 8496 1619 8512
rect 219 8450 1619 8466
rect 219 8416 231 8450
rect 1607 8416 1619 8450
rect 219 8400 1619 8416
rect 219 8354 1619 8370
rect 219 8320 231 8354
rect 1607 8320 1619 8354
rect 219 8304 1619 8320
rect 219 8258 1619 8274
rect 219 8224 231 8258
rect 1607 8224 1619 8258
rect 219 8208 1619 8224
rect 219 8162 1619 8178
rect 219 8128 231 8162
rect 1607 8128 1619 8162
rect 219 8112 1619 8128
rect 219 8066 1619 8082
rect 219 8032 231 8066
rect 1607 8032 1619 8066
rect 219 8016 1619 8032
rect 219 7970 1619 7986
rect 219 7936 231 7970
rect 1607 7936 1619 7970
rect 219 7920 1619 7936
rect 219 7874 1619 7890
rect 219 7840 231 7874
rect 1607 7840 1619 7874
rect 219 7824 1619 7840
rect 219 7778 1619 7794
rect 219 7744 231 7778
rect 1607 7744 1619 7778
rect 219 7728 1619 7744
rect 219 7682 1619 7698
rect 219 7648 231 7682
rect 1607 7648 1619 7682
rect 219 7632 1619 7648
rect 219 7586 1619 7602
rect 219 7552 231 7586
rect 1607 7552 1619 7586
rect 219 7536 1619 7552
rect 219 7490 1619 7506
rect 219 7456 231 7490
rect 1607 7456 1619 7490
rect 219 7440 1619 7456
rect 219 7394 1619 7410
rect 219 7360 231 7394
rect 1607 7360 1619 7394
rect 219 7344 1619 7360
rect 219 7298 1619 7314
rect 219 7264 231 7298
rect 1607 7264 1619 7298
rect 219 7248 1619 7264
rect 219 7202 1619 7218
rect 219 7168 231 7202
rect 1607 7168 1619 7202
rect 219 7152 1619 7168
rect 219 7106 1619 7122
rect 219 7072 231 7106
rect 1607 7072 1619 7106
rect 219 7056 1619 7072
rect 219 7010 1619 7026
rect 219 6976 231 7010
rect 1607 6976 1619 7010
rect 219 6960 1619 6976
rect 219 6914 1619 6930
rect 219 6880 231 6914
rect 1607 6880 1619 6914
rect 219 6864 1619 6880
rect 219 6818 1619 6834
rect 219 6784 231 6818
rect 1607 6784 1619 6818
rect 219 6768 1619 6784
rect 219 6722 1619 6738
rect 219 6688 231 6722
rect 1607 6688 1619 6722
rect 219 6672 1619 6688
rect 219 6626 1619 6642
rect 219 6592 231 6626
rect 1607 6592 1619 6626
rect 219 6576 1619 6592
rect 219 6530 1619 6546
rect 219 6496 231 6530
rect 1607 6496 1619 6530
rect 219 6480 1619 6496
rect 219 6434 1619 6450
rect 219 6400 231 6434
rect 1607 6400 1619 6434
rect 219 6384 1619 6400
rect 219 6338 1619 6354
rect 219 6304 231 6338
rect 1607 6304 1619 6338
rect 219 6288 1619 6304
rect 219 6242 1619 6258
rect 219 6208 231 6242
rect 1607 6208 1619 6242
rect 219 6192 1619 6208
rect 219 6146 1619 6162
rect 219 6112 231 6146
rect 1607 6112 1619 6146
rect 219 6096 1619 6112
rect 219 6050 1619 6066
rect 219 6016 231 6050
rect 1607 6016 1619 6050
rect 219 6000 1619 6016
rect 219 5954 1619 5970
rect 219 5920 231 5954
rect 1607 5920 1619 5954
rect 219 5904 1619 5920
rect 219 5858 1619 5874
rect 219 5824 231 5858
rect 1607 5824 1619 5858
rect 219 5808 1619 5824
rect 219 5762 1619 5778
rect 219 5728 231 5762
rect 1607 5728 1619 5762
rect 219 5712 1619 5728
rect 219 5666 1619 5682
rect 219 5632 231 5666
rect 1607 5632 1619 5666
rect 219 5616 1619 5632
rect 219 5570 1619 5586
rect 219 5536 231 5570
rect 1607 5536 1619 5570
rect 219 5520 1619 5536
rect 219 5474 1619 5490
rect 219 5440 231 5474
rect 1607 5440 1619 5474
rect 219 5424 1619 5440
rect 219 5378 1619 5394
rect 219 5344 231 5378
rect 1607 5344 1619 5378
rect 219 5328 1619 5344
rect 219 5282 1619 5298
rect 219 5248 231 5282
rect 1607 5248 1619 5282
rect 219 5232 1619 5248
rect 219 5186 1619 5202
rect 219 5152 231 5186
rect 1607 5152 1619 5186
rect 219 5136 1619 5152
rect 219 5090 1619 5106
rect 219 5056 231 5090
rect 1607 5056 1619 5090
rect 219 5040 1619 5056
rect 219 4994 1619 5010
rect 219 4960 231 4994
rect 1607 4960 1619 4994
rect 219 4944 1619 4960
rect 219 4898 1619 4914
rect 219 4864 231 4898
rect 1607 4864 1619 4898
rect 219 4848 1619 4864
rect 219 4802 1619 4818
rect 219 4768 231 4802
rect 1607 4768 1619 4802
rect 219 4752 1619 4768
rect 219 4706 1619 4722
rect 219 4672 231 4706
rect 1607 4672 1619 4706
rect 219 4656 1619 4672
rect 219 4610 1619 4626
rect 219 4576 231 4610
rect 1607 4576 1619 4610
rect 219 4560 1619 4576
rect 219 4514 1619 4530
rect 219 4480 231 4514
rect 1607 4480 1619 4514
rect 219 4464 1619 4480
rect 219 4418 1619 4434
rect 219 4384 231 4418
rect 1607 4384 1619 4418
rect 219 4368 1619 4384
rect 219 4322 1619 4338
rect 219 4288 231 4322
rect 1607 4288 1619 4322
rect 219 4272 1619 4288
rect 219 4226 1619 4242
rect 219 4192 231 4226
rect 1607 4192 1619 4226
rect 219 4176 1619 4192
rect 219 4130 1619 4146
rect 219 4096 231 4130
rect 1607 4096 1619 4130
rect 219 4080 1619 4096
rect 219 4034 1619 4050
rect 219 4000 231 4034
rect 1607 4000 1619 4034
rect 219 3984 1619 4000
rect 219 3938 1619 3954
rect 219 3904 231 3938
rect 1607 3904 1619 3938
rect 219 3888 1619 3904
rect 219 3842 1619 3858
rect 219 3808 231 3842
rect 1607 3808 1619 3842
rect 219 3792 1619 3808
rect 219 3746 1619 3762
rect 219 3712 231 3746
rect 1607 3712 1619 3746
rect 219 3696 1619 3712
rect 219 3650 1619 3666
rect 219 3616 231 3650
rect 1607 3616 1619 3650
rect 219 3600 1619 3616
rect 219 3554 1619 3570
rect 219 3520 231 3554
rect 1607 3520 1619 3554
rect 219 3504 1619 3520
rect 219 3458 1619 3474
rect 219 3424 231 3458
rect 1607 3424 1619 3458
rect 219 3408 1619 3424
rect 219 3362 1619 3378
rect 219 3328 231 3362
rect 1607 3328 1619 3362
rect 219 3312 1619 3328
rect 219 3266 1619 3282
rect 219 3232 231 3266
rect 1607 3232 1619 3266
rect 219 3216 1619 3232
rect 219 3170 1619 3186
rect 219 3136 231 3170
rect 1607 3136 1619 3170
rect 219 3120 1619 3136
rect 219 3074 1619 3090
rect 219 3040 231 3074
rect 1607 3040 1619 3074
rect 219 3024 1619 3040
rect 219 2978 1619 2994
rect 219 2944 231 2978
rect 1607 2944 1619 2978
rect 219 2928 1619 2944
rect 219 2882 1619 2898
rect 219 2848 231 2882
rect 1607 2848 1619 2882
rect 219 2832 1619 2848
rect 219 2786 1619 2802
rect 219 2752 231 2786
rect 1607 2752 1619 2786
rect 219 2736 1619 2752
rect 219 2690 1619 2706
rect 219 2656 231 2690
rect 1607 2656 1619 2690
rect 219 2640 1619 2656
rect 219 2594 1619 2610
rect 219 2560 231 2594
rect 1607 2560 1619 2594
rect 219 2544 1619 2560
rect 219 2498 1619 2514
rect 219 2464 231 2498
rect 1607 2464 1619 2498
rect 219 2448 1619 2464
rect 219 2402 1619 2418
rect 219 2368 231 2402
rect 1607 2368 1619 2402
rect 219 2352 1619 2368
rect 219 2306 1619 2322
rect 219 2272 231 2306
rect 1607 2272 1619 2306
rect 219 2256 1619 2272
rect 219 2210 1619 2226
rect 219 2176 231 2210
rect 1607 2176 1619 2210
rect 219 2160 1619 2176
rect 219 2114 1619 2130
rect 219 2080 231 2114
rect 1607 2080 1619 2114
rect 219 2064 1619 2080
rect 219 2018 1619 2034
rect 219 1984 231 2018
rect 1607 1984 1619 2018
rect 219 1968 1619 1984
rect 219 1922 1619 1938
rect 219 1888 231 1922
rect 1607 1888 1619 1922
rect 219 1872 1619 1888
rect 219 1826 1619 1842
rect 219 1792 231 1826
rect 1607 1792 1619 1826
rect 219 1776 1619 1792
rect 219 1730 1619 1746
rect 219 1696 231 1730
rect 1607 1696 1619 1730
rect 219 1680 1619 1696
rect 219 1634 1619 1650
rect 219 1600 231 1634
rect 1607 1600 1619 1634
rect 219 1584 1619 1600
rect 219 1538 1619 1554
rect 219 1504 231 1538
rect 1607 1504 1619 1538
rect 219 1488 1619 1504
rect 219 1442 1619 1458
rect 219 1408 231 1442
rect 1607 1408 1619 1442
rect 219 1392 1619 1408
rect 219 1346 1619 1362
rect 219 1312 231 1346
rect 1607 1312 1619 1346
rect 219 1296 1619 1312
rect 219 1250 1619 1266
rect 219 1216 231 1250
rect 1607 1216 1619 1250
rect 219 1200 1619 1216
rect 219 1154 1619 1170
rect 219 1120 231 1154
rect 1607 1120 1619 1154
rect 219 1104 1619 1120
rect 219 1058 1619 1074
rect 219 1024 231 1058
rect 1607 1024 1619 1058
rect 219 1008 1619 1024
rect 219 962 1619 978
rect 219 928 231 962
rect 1607 928 1619 962
rect 219 912 1619 928
rect 219 866 1619 882
rect 219 832 231 866
rect 1607 832 1619 866
rect 219 816 1619 832
rect 219 770 1619 786
rect 219 736 231 770
rect 1607 736 1619 770
rect 219 720 1619 736
rect 219 674 1619 690
rect 219 640 231 674
rect 1607 640 1619 674
rect 219 628 1619 640
<< pdiffc >>
rect 231 21760 1607 21794
rect 231 21664 1607 21698
rect 231 21568 1607 21602
rect 231 21472 1607 21506
rect 231 21376 1607 21410
rect 231 21280 1607 21314
rect 231 21184 1607 21218
rect 231 21088 1607 21122
rect 231 20992 1607 21026
rect 231 20896 1607 20930
rect 231 20800 1607 20834
rect 231 20704 1607 20738
rect 231 20608 1607 20642
rect 231 20512 1607 20546
rect 231 20416 1607 20450
rect 231 20320 1607 20354
rect 231 20224 1607 20258
rect 231 20128 1607 20162
rect 231 20032 1607 20066
rect 231 19936 1607 19970
rect 231 19840 1607 19874
rect 231 19744 1607 19778
rect 231 19648 1607 19682
rect 231 19552 1607 19586
rect 231 19456 1607 19490
rect 231 19360 1607 19394
rect 231 19264 1607 19298
rect 231 19168 1607 19202
rect 231 19072 1607 19106
rect 231 18976 1607 19010
rect 231 18880 1607 18914
rect 231 18784 1607 18818
rect 231 18688 1607 18722
rect 231 18592 1607 18626
rect 231 18496 1607 18530
rect 231 18400 1607 18434
rect 231 18304 1607 18338
rect 231 18208 1607 18242
rect 231 18112 1607 18146
rect 231 18016 1607 18050
rect 231 17920 1607 17954
rect 231 17824 1607 17858
rect 231 17728 1607 17762
rect 231 17632 1607 17666
rect 231 17536 1607 17570
rect 231 17440 1607 17474
rect 231 17344 1607 17378
rect 231 17248 1607 17282
rect 231 17152 1607 17186
rect 231 17056 1607 17090
rect 231 16960 1607 16994
rect 231 16864 1607 16898
rect 231 16768 1607 16802
rect 231 16672 1607 16706
rect 231 16576 1607 16610
rect 231 16480 1607 16514
rect 231 16384 1607 16418
rect 231 16288 1607 16322
rect 231 16192 1607 16226
rect 231 16096 1607 16130
rect 231 16000 1607 16034
rect 231 15904 1607 15938
rect 231 15808 1607 15842
rect 231 15712 1607 15746
rect 231 15616 1607 15650
rect 231 15520 1607 15554
rect 231 15424 1607 15458
rect 231 15328 1607 15362
rect 231 15232 1607 15266
rect 231 15136 1607 15170
rect 231 15040 1607 15074
rect 231 14944 1607 14978
rect 231 14848 1607 14882
rect 231 14752 1607 14786
rect 231 14656 1607 14690
rect 231 14560 1607 14594
rect 231 14464 1607 14498
rect 231 14368 1607 14402
rect 231 14272 1607 14306
rect 231 14176 1607 14210
rect 231 14080 1607 14114
rect 231 13984 1607 14018
rect 231 13888 1607 13922
rect 231 13792 1607 13826
rect 231 13696 1607 13730
rect 231 13600 1607 13634
rect 231 13504 1607 13538
rect 231 13408 1607 13442
rect 231 13312 1607 13346
rect 231 13216 1607 13250
rect 231 13120 1607 13154
rect 231 13024 1607 13058
rect 231 12928 1607 12962
rect 231 12832 1607 12866
rect 231 12736 1607 12770
rect 231 12640 1607 12674
rect 231 12544 1607 12578
rect 231 12448 1607 12482
rect 231 12352 1607 12386
rect 231 12256 1607 12290
rect 231 12160 1607 12194
rect 231 12064 1607 12098
rect 231 11968 1607 12002
rect 231 11872 1607 11906
rect 231 11776 1607 11810
rect 231 11680 1607 11714
rect 231 11584 1607 11618
rect 231 11488 1607 11522
rect 231 11392 1607 11426
rect 231 11296 1607 11330
rect 231 11200 1607 11234
rect 231 11104 1607 11138
rect 231 11008 1607 11042
rect 231 10912 1607 10946
rect 231 10816 1607 10850
rect 231 10720 1607 10754
rect 231 10624 1607 10658
rect 231 10528 1607 10562
rect 231 10432 1607 10466
rect 231 10336 1607 10370
rect 231 10240 1607 10274
rect 231 10144 1607 10178
rect 231 10048 1607 10082
rect 231 9952 1607 9986
rect 231 9856 1607 9890
rect 231 9760 1607 9794
rect 231 9664 1607 9698
rect 231 9568 1607 9602
rect 231 9472 1607 9506
rect 231 9376 1607 9410
rect 231 9280 1607 9314
rect 231 9184 1607 9218
rect 231 9088 1607 9122
rect 231 8992 1607 9026
rect 231 8896 1607 8930
rect 231 8800 1607 8834
rect 231 8704 1607 8738
rect 231 8608 1607 8642
rect 231 8512 1607 8546
rect 231 8416 1607 8450
rect 231 8320 1607 8354
rect 231 8224 1607 8258
rect 231 8128 1607 8162
rect 231 8032 1607 8066
rect 231 7936 1607 7970
rect 231 7840 1607 7874
rect 231 7744 1607 7778
rect 231 7648 1607 7682
rect 231 7552 1607 7586
rect 231 7456 1607 7490
rect 231 7360 1607 7394
rect 231 7264 1607 7298
rect 231 7168 1607 7202
rect 231 7072 1607 7106
rect 231 6976 1607 7010
rect 231 6880 1607 6914
rect 231 6784 1607 6818
rect 231 6688 1607 6722
rect 231 6592 1607 6626
rect 231 6496 1607 6530
rect 231 6400 1607 6434
rect 231 6304 1607 6338
rect 231 6208 1607 6242
rect 231 6112 1607 6146
rect 231 6016 1607 6050
rect 231 5920 1607 5954
rect 231 5824 1607 5858
rect 231 5728 1607 5762
rect 231 5632 1607 5666
rect 231 5536 1607 5570
rect 231 5440 1607 5474
rect 231 5344 1607 5378
rect 231 5248 1607 5282
rect 231 5152 1607 5186
rect 231 5056 1607 5090
rect 231 4960 1607 4994
rect 231 4864 1607 4898
rect 231 4768 1607 4802
rect 231 4672 1607 4706
rect 231 4576 1607 4610
rect 231 4480 1607 4514
rect 231 4384 1607 4418
rect 231 4288 1607 4322
rect 231 4192 1607 4226
rect 231 4096 1607 4130
rect 231 4000 1607 4034
rect 231 3904 1607 3938
rect 231 3808 1607 3842
rect 231 3712 1607 3746
rect 231 3616 1607 3650
rect 231 3520 1607 3554
rect 231 3424 1607 3458
rect 231 3328 1607 3362
rect 231 3232 1607 3266
rect 231 3136 1607 3170
rect 231 3040 1607 3074
rect 231 2944 1607 2978
rect 231 2848 1607 2882
rect 231 2752 1607 2786
rect 231 2656 1607 2690
rect 231 2560 1607 2594
rect 231 2464 1607 2498
rect 231 2368 1607 2402
rect 231 2272 1607 2306
rect 231 2176 1607 2210
rect 231 2080 1607 2114
rect 231 1984 1607 2018
rect 231 1888 1607 1922
rect 231 1792 1607 1826
rect 231 1696 1607 1730
rect 231 1600 1607 1634
rect 231 1504 1607 1538
rect 231 1408 1607 1442
rect 231 1312 1607 1346
rect 231 1216 1607 1250
rect 231 1120 1607 1154
rect 231 1024 1607 1058
rect 231 928 1607 962
rect 231 832 1607 866
rect 231 736 1607 770
rect 231 640 1607 674
<< nsubdiff >>
rect 36 21874 132 21908
rect 1706 21874 1802 21908
rect 36 21812 70 21874
rect 1768 21812 1802 21874
rect 36 560 70 622
rect 1768 560 1802 622
rect 36 526 132 560
rect 1706 526 1802 560
<< nsubdiffcont >>
rect 132 21874 1706 21908
rect 36 622 70 21812
rect 1768 622 1802 21812
rect 132 526 1706 560
<< poly >>
rect 122 21746 188 21762
rect 122 21712 138 21746
rect 172 21744 188 21746
rect 172 21714 219 21744
rect 1619 21714 1645 21744
rect 172 21712 188 21714
rect 122 21696 188 21712
rect 1650 21650 1716 21666
rect 1650 21648 1666 21650
rect 193 21618 219 21648
rect 1619 21618 1666 21648
rect 122 21554 188 21570
rect 122 21520 138 21554
rect 172 21552 188 21554
rect 1650 21616 1666 21618
rect 1700 21616 1716 21650
rect 1650 21600 1716 21616
rect 172 21522 219 21552
rect 1619 21522 1645 21552
rect 172 21520 188 21522
rect 122 21504 188 21520
rect 1650 21458 1716 21474
rect 1650 21456 1666 21458
rect 193 21426 219 21456
rect 1619 21426 1666 21456
rect 122 21362 188 21378
rect 122 21328 138 21362
rect 172 21360 188 21362
rect 1650 21424 1666 21426
rect 1700 21424 1716 21458
rect 1650 21408 1716 21424
rect 172 21330 219 21360
rect 1619 21330 1645 21360
rect 172 21328 188 21330
rect 122 21312 188 21328
rect 1650 21266 1716 21282
rect 1650 21264 1666 21266
rect 193 21234 219 21264
rect 1619 21234 1666 21264
rect 122 21170 188 21186
rect 122 21136 138 21170
rect 172 21168 188 21170
rect 1650 21232 1666 21234
rect 1700 21232 1716 21266
rect 1650 21216 1716 21232
rect 172 21138 219 21168
rect 1619 21138 1645 21168
rect 172 21136 188 21138
rect 122 21120 188 21136
rect 1650 21074 1716 21090
rect 1650 21072 1666 21074
rect 193 21042 219 21072
rect 1619 21042 1666 21072
rect 122 20978 188 20994
rect 122 20944 138 20978
rect 172 20976 188 20978
rect 1650 21040 1666 21042
rect 1700 21040 1716 21074
rect 1650 21024 1716 21040
rect 172 20946 219 20976
rect 1619 20946 1645 20976
rect 172 20944 188 20946
rect 122 20928 188 20944
rect 1650 20882 1716 20898
rect 1650 20880 1666 20882
rect 193 20850 219 20880
rect 1619 20850 1666 20880
rect 122 20786 188 20802
rect 122 20752 138 20786
rect 172 20784 188 20786
rect 1650 20848 1666 20850
rect 1700 20848 1716 20882
rect 1650 20832 1716 20848
rect 172 20754 219 20784
rect 1619 20754 1645 20784
rect 172 20752 188 20754
rect 122 20736 188 20752
rect 1650 20690 1716 20706
rect 1650 20688 1666 20690
rect 193 20658 219 20688
rect 1619 20658 1666 20688
rect 122 20594 188 20610
rect 122 20560 138 20594
rect 172 20592 188 20594
rect 1650 20656 1666 20658
rect 1700 20656 1716 20690
rect 1650 20640 1716 20656
rect 172 20562 219 20592
rect 1619 20562 1645 20592
rect 172 20560 188 20562
rect 122 20544 188 20560
rect 1650 20498 1716 20514
rect 1650 20496 1666 20498
rect 193 20466 219 20496
rect 1619 20466 1666 20496
rect 122 20402 188 20418
rect 122 20368 138 20402
rect 172 20400 188 20402
rect 1650 20464 1666 20466
rect 1700 20464 1716 20498
rect 1650 20448 1716 20464
rect 172 20370 219 20400
rect 1619 20370 1645 20400
rect 172 20368 188 20370
rect 122 20352 188 20368
rect 1650 20306 1716 20322
rect 1650 20304 1666 20306
rect 193 20274 219 20304
rect 1619 20274 1666 20304
rect 122 20210 188 20226
rect 122 20176 138 20210
rect 172 20208 188 20210
rect 1650 20272 1666 20274
rect 1700 20272 1716 20306
rect 1650 20256 1716 20272
rect 172 20178 219 20208
rect 1619 20178 1645 20208
rect 172 20176 188 20178
rect 122 20160 188 20176
rect 1650 20114 1716 20130
rect 1650 20112 1666 20114
rect 193 20082 219 20112
rect 1619 20082 1666 20112
rect 122 20018 188 20034
rect 122 19984 138 20018
rect 172 20016 188 20018
rect 1650 20080 1666 20082
rect 1700 20080 1716 20114
rect 1650 20064 1716 20080
rect 172 19986 219 20016
rect 1619 19986 1645 20016
rect 172 19984 188 19986
rect 122 19968 188 19984
rect 1650 19922 1716 19938
rect 1650 19920 1666 19922
rect 193 19890 219 19920
rect 1619 19890 1666 19920
rect 122 19826 188 19842
rect 122 19792 138 19826
rect 172 19824 188 19826
rect 1650 19888 1666 19890
rect 1700 19888 1716 19922
rect 1650 19872 1716 19888
rect 172 19794 219 19824
rect 1619 19794 1645 19824
rect 172 19792 188 19794
rect 122 19776 188 19792
rect 1650 19730 1716 19746
rect 1650 19728 1666 19730
rect 193 19698 219 19728
rect 1619 19698 1666 19728
rect 122 19634 188 19650
rect 122 19600 138 19634
rect 172 19632 188 19634
rect 1650 19696 1666 19698
rect 1700 19696 1716 19730
rect 1650 19680 1716 19696
rect 172 19602 219 19632
rect 1619 19602 1645 19632
rect 172 19600 188 19602
rect 122 19584 188 19600
rect 1650 19538 1716 19554
rect 1650 19536 1666 19538
rect 193 19506 219 19536
rect 1619 19506 1666 19536
rect 122 19442 188 19458
rect 122 19408 138 19442
rect 172 19440 188 19442
rect 1650 19504 1666 19506
rect 1700 19504 1716 19538
rect 1650 19488 1716 19504
rect 172 19410 219 19440
rect 1619 19410 1645 19440
rect 172 19408 188 19410
rect 122 19392 188 19408
rect 1650 19346 1716 19362
rect 1650 19344 1666 19346
rect 193 19314 219 19344
rect 1619 19314 1666 19344
rect 122 19250 188 19266
rect 122 19216 138 19250
rect 172 19248 188 19250
rect 1650 19312 1666 19314
rect 1700 19312 1716 19346
rect 1650 19296 1716 19312
rect 172 19218 219 19248
rect 1619 19218 1645 19248
rect 172 19216 188 19218
rect 122 19200 188 19216
rect 1650 19154 1716 19170
rect 1650 19152 1666 19154
rect 193 19122 219 19152
rect 1619 19122 1666 19152
rect 122 19058 188 19074
rect 122 19024 138 19058
rect 172 19056 188 19058
rect 1650 19120 1666 19122
rect 1700 19120 1716 19154
rect 1650 19104 1716 19120
rect 172 19026 219 19056
rect 1619 19026 1645 19056
rect 172 19024 188 19026
rect 122 19008 188 19024
rect 1650 18962 1716 18978
rect 1650 18960 1666 18962
rect 193 18930 219 18960
rect 1619 18930 1666 18960
rect 122 18866 188 18882
rect 122 18832 138 18866
rect 172 18864 188 18866
rect 1650 18928 1666 18930
rect 1700 18928 1716 18962
rect 1650 18912 1716 18928
rect 172 18834 219 18864
rect 1619 18834 1645 18864
rect 172 18832 188 18834
rect 122 18816 188 18832
rect 1650 18770 1716 18786
rect 1650 18768 1666 18770
rect 193 18738 219 18768
rect 1619 18738 1666 18768
rect 122 18674 188 18690
rect 122 18640 138 18674
rect 172 18672 188 18674
rect 1650 18736 1666 18738
rect 1700 18736 1716 18770
rect 1650 18720 1716 18736
rect 172 18642 219 18672
rect 1619 18642 1645 18672
rect 172 18640 188 18642
rect 122 18624 188 18640
rect 1650 18578 1716 18594
rect 1650 18576 1666 18578
rect 193 18546 219 18576
rect 1619 18546 1666 18576
rect 122 18482 188 18498
rect 122 18448 138 18482
rect 172 18480 188 18482
rect 1650 18544 1666 18546
rect 1700 18544 1716 18578
rect 1650 18528 1716 18544
rect 172 18450 219 18480
rect 1619 18450 1645 18480
rect 172 18448 188 18450
rect 122 18432 188 18448
rect 1650 18386 1716 18402
rect 1650 18384 1666 18386
rect 193 18354 219 18384
rect 1619 18354 1666 18384
rect 122 18290 188 18306
rect 122 18256 138 18290
rect 172 18288 188 18290
rect 1650 18352 1666 18354
rect 1700 18352 1716 18386
rect 1650 18336 1716 18352
rect 172 18258 219 18288
rect 1619 18258 1645 18288
rect 172 18256 188 18258
rect 122 18240 188 18256
rect 1650 18194 1716 18210
rect 1650 18192 1666 18194
rect 193 18162 219 18192
rect 1619 18162 1666 18192
rect 122 18098 188 18114
rect 122 18064 138 18098
rect 172 18096 188 18098
rect 1650 18160 1666 18162
rect 1700 18160 1716 18194
rect 1650 18144 1716 18160
rect 172 18066 219 18096
rect 1619 18066 1645 18096
rect 172 18064 188 18066
rect 122 18048 188 18064
rect 1650 18002 1716 18018
rect 1650 18000 1666 18002
rect 193 17970 219 18000
rect 1619 17970 1666 18000
rect 122 17906 188 17922
rect 122 17872 138 17906
rect 172 17904 188 17906
rect 1650 17968 1666 17970
rect 1700 17968 1716 18002
rect 1650 17952 1716 17968
rect 172 17874 219 17904
rect 1619 17874 1645 17904
rect 172 17872 188 17874
rect 122 17856 188 17872
rect 1650 17810 1716 17826
rect 1650 17808 1666 17810
rect 193 17778 219 17808
rect 1619 17778 1666 17808
rect 122 17714 188 17730
rect 122 17680 138 17714
rect 172 17712 188 17714
rect 1650 17776 1666 17778
rect 1700 17776 1716 17810
rect 1650 17760 1716 17776
rect 172 17682 219 17712
rect 1619 17682 1645 17712
rect 172 17680 188 17682
rect 122 17664 188 17680
rect 1650 17618 1716 17634
rect 1650 17616 1666 17618
rect 193 17586 219 17616
rect 1619 17586 1666 17616
rect 122 17522 188 17538
rect 122 17488 138 17522
rect 172 17520 188 17522
rect 1650 17584 1666 17586
rect 1700 17584 1716 17618
rect 1650 17568 1716 17584
rect 172 17490 219 17520
rect 1619 17490 1645 17520
rect 172 17488 188 17490
rect 122 17472 188 17488
rect 1650 17426 1716 17442
rect 1650 17424 1666 17426
rect 193 17394 219 17424
rect 1619 17394 1666 17424
rect 122 17330 188 17346
rect 122 17296 138 17330
rect 172 17328 188 17330
rect 1650 17392 1666 17394
rect 1700 17392 1716 17426
rect 1650 17376 1716 17392
rect 172 17298 219 17328
rect 1619 17298 1645 17328
rect 172 17296 188 17298
rect 122 17280 188 17296
rect 1650 17234 1716 17250
rect 1650 17232 1666 17234
rect 193 17202 219 17232
rect 1619 17202 1666 17232
rect 122 17138 188 17154
rect 122 17104 138 17138
rect 172 17136 188 17138
rect 1650 17200 1666 17202
rect 1700 17200 1716 17234
rect 1650 17184 1716 17200
rect 172 17106 219 17136
rect 1619 17106 1645 17136
rect 172 17104 188 17106
rect 122 17088 188 17104
rect 1650 17042 1716 17058
rect 1650 17040 1666 17042
rect 193 17010 219 17040
rect 1619 17010 1666 17040
rect 122 16946 188 16962
rect 122 16912 138 16946
rect 172 16944 188 16946
rect 1650 17008 1666 17010
rect 1700 17008 1716 17042
rect 1650 16992 1716 17008
rect 172 16914 219 16944
rect 1619 16914 1645 16944
rect 172 16912 188 16914
rect 122 16896 188 16912
rect 1650 16850 1716 16866
rect 1650 16848 1666 16850
rect 193 16818 219 16848
rect 1619 16818 1666 16848
rect 122 16754 188 16770
rect 122 16720 138 16754
rect 172 16752 188 16754
rect 1650 16816 1666 16818
rect 1700 16816 1716 16850
rect 1650 16800 1716 16816
rect 172 16722 219 16752
rect 1619 16722 1645 16752
rect 172 16720 188 16722
rect 122 16704 188 16720
rect 1650 16658 1716 16674
rect 1650 16656 1666 16658
rect 193 16626 219 16656
rect 1619 16626 1666 16656
rect 122 16562 188 16578
rect 122 16528 138 16562
rect 172 16560 188 16562
rect 1650 16624 1666 16626
rect 1700 16624 1716 16658
rect 1650 16608 1716 16624
rect 172 16530 219 16560
rect 1619 16530 1645 16560
rect 172 16528 188 16530
rect 122 16512 188 16528
rect 1650 16466 1716 16482
rect 1650 16464 1666 16466
rect 193 16434 219 16464
rect 1619 16434 1666 16464
rect 122 16370 188 16386
rect 122 16336 138 16370
rect 172 16368 188 16370
rect 1650 16432 1666 16434
rect 1700 16432 1716 16466
rect 1650 16416 1716 16432
rect 172 16338 219 16368
rect 1619 16338 1645 16368
rect 172 16336 188 16338
rect 122 16320 188 16336
rect 1650 16274 1716 16290
rect 1650 16272 1666 16274
rect 193 16242 219 16272
rect 1619 16242 1666 16272
rect 122 16178 188 16194
rect 122 16144 138 16178
rect 172 16176 188 16178
rect 1650 16240 1666 16242
rect 1700 16240 1716 16274
rect 1650 16224 1716 16240
rect 172 16146 219 16176
rect 1619 16146 1645 16176
rect 172 16144 188 16146
rect 122 16128 188 16144
rect 1650 16082 1716 16098
rect 1650 16080 1666 16082
rect 193 16050 219 16080
rect 1619 16050 1666 16080
rect 122 15986 188 16002
rect 122 15952 138 15986
rect 172 15984 188 15986
rect 1650 16048 1666 16050
rect 1700 16048 1716 16082
rect 1650 16032 1716 16048
rect 172 15954 219 15984
rect 1619 15954 1645 15984
rect 172 15952 188 15954
rect 122 15936 188 15952
rect 1650 15890 1716 15906
rect 1650 15888 1666 15890
rect 193 15858 219 15888
rect 1619 15858 1666 15888
rect 122 15794 188 15810
rect 122 15760 138 15794
rect 172 15792 188 15794
rect 1650 15856 1666 15858
rect 1700 15856 1716 15890
rect 1650 15840 1716 15856
rect 172 15762 219 15792
rect 1619 15762 1645 15792
rect 172 15760 188 15762
rect 122 15744 188 15760
rect 1650 15698 1716 15714
rect 1650 15696 1666 15698
rect 193 15666 219 15696
rect 1619 15666 1666 15696
rect 122 15602 188 15618
rect 122 15568 138 15602
rect 172 15600 188 15602
rect 1650 15664 1666 15666
rect 1700 15664 1716 15698
rect 1650 15648 1716 15664
rect 172 15570 219 15600
rect 1619 15570 1645 15600
rect 172 15568 188 15570
rect 122 15552 188 15568
rect 1650 15506 1716 15522
rect 1650 15504 1666 15506
rect 193 15474 219 15504
rect 1619 15474 1666 15504
rect 122 15410 188 15426
rect 122 15376 138 15410
rect 172 15408 188 15410
rect 1650 15472 1666 15474
rect 1700 15472 1716 15506
rect 1650 15456 1716 15472
rect 172 15378 219 15408
rect 1619 15378 1645 15408
rect 172 15376 188 15378
rect 122 15360 188 15376
rect 1650 15314 1716 15330
rect 1650 15312 1666 15314
rect 193 15282 219 15312
rect 1619 15282 1666 15312
rect 122 15218 188 15234
rect 122 15184 138 15218
rect 172 15216 188 15218
rect 1650 15280 1666 15282
rect 1700 15280 1716 15314
rect 1650 15264 1716 15280
rect 172 15186 219 15216
rect 1619 15186 1645 15216
rect 172 15184 188 15186
rect 122 15168 188 15184
rect 1650 15122 1716 15138
rect 1650 15120 1666 15122
rect 193 15090 219 15120
rect 1619 15090 1666 15120
rect 122 15026 188 15042
rect 122 14992 138 15026
rect 172 15024 188 15026
rect 1650 15088 1666 15090
rect 1700 15088 1716 15122
rect 1650 15072 1716 15088
rect 172 14994 219 15024
rect 1619 14994 1645 15024
rect 172 14992 188 14994
rect 122 14976 188 14992
rect 1650 14930 1716 14946
rect 1650 14928 1666 14930
rect 193 14898 219 14928
rect 1619 14898 1666 14928
rect 122 14834 188 14850
rect 122 14800 138 14834
rect 172 14832 188 14834
rect 1650 14896 1666 14898
rect 1700 14896 1716 14930
rect 1650 14880 1716 14896
rect 172 14802 219 14832
rect 1619 14802 1645 14832
rect 172 14800 188 14802
rect 122 14784 188 14800
rect 1650 14738 1716 14754
rect 1650 14736 1666 14738
rect 193 14706 219 14736
rect 1619 14706 1666 14736
rect 122 14642 188 14658
rect 122 14608 138 14642
rect 172 14640 188 14642
rect 1650 14704 1666 14706
rect 1700 14704 1716 14738
rect 1650 14688 1716 14704
rect 172 14610 219 14640
rect 1619 14610 1645 14640
rect 172 14608 188 14610
rect 122 14592 188 14608
rect 1650 14546 1716 14562
rect 1650 14544 1666 14546
rect 193 14514 219 14544
rect 1619 14514 1666 14544
rect 122 14450 188 14466
rect 122 14416 138 14450
rect 172 14448 188 14450
rect 1650 14512 1666 14514
rect 1700 14512 1716 14546
rect 1650 14496 1716 14512
rect 172 14418 219 14448
rect 1619 14418 1645 14448
rect 172 14416 188 14418
rect 122 14400 188 14416
rect 1650 14354 1716 14370
rect 1650 14352 1666 14354
rect 193 14322 219 14352
rect 1619 14322 1666 14352
rect 122 14258 188 14274
rect 122 14224 138 14258
rect 172 14256 188 14258
rect 1650 14320 1666 14322
rect 1700 14320 1716 14354
rect 1650 14304 1716 14320
rect 172 14226 219 14256
rect 1619 14226 1645 14256
rect 172 14224 188 14226
rect 122 14208 188 14224
rect 1650 14162 1716 14178
rect 1650 14160 1666 14162
rect 193 14130 219 14160
rect 1619 14130 1666 14160
rect 122 14066 188 14082
rect 122 14032 138 14066
rect 172 14064 188 14066
rect 1650 14128 1666 14130
rect 1700 14128 1716 14162
rect 1650 14112 1716 14128
rect 172 14034 219 14064
rect 1619 14034 1645 14064
rect 172 14032 188 14034
rect 122 14016 188 14032
rect 1650 13970 1716 13986
rect 1650 13968 1666 13970
rect 193 13938 219 13968
rect 1619 13938 1666 13968
rect 122 13874 188 13890
rect 122 13840 138 13874
rect 172 13872 188 13874
rect 1650 13936 1666 13938
rect 1700 13936 1716 13970
rect 1650 13920 1716 13936
rect 172 13842 219 13872
rect 1619 13842 1645 13872
rect 172 13840 188 13842
rect 122 13824 188 13840
rect 1650 13778 1716 13794
rect 1650 13776 1666 13778
rect 193 13746 219 13776
rect 1619 13746 1666 13776
rect 122 13682 188 13698
rect 122 13648 138 13682
rect 172 13680 188 13682
rect 1650 13744 1666 13746
rect 1700 13744 1716 13778
rect 1650 13728 1716 13744
rect 172 13650 219 13680
rect 1619 13650 1645 13680
rect 172 13648 188 13650
rect 122 13632 188 13648
rect 1650 13586 1716 13602
rect 1650 13584 1666 13586
rect 193 13554 219 13584
rect 1619 13554 1666 13584
rect 122 13490 188 13506
rect 122 13456 138 13490
rect 172 13488 188 13490
rect 1650 13552 1666 13554
rect 1700 13552 1716 13586
rect 1650 13536 1716 13552
rect 172 13458 219 13488
rect 1619 13458 1645 13488
rect 172 13456 188 13458
rect 122 13440 188 13456
rect 1650 13394 1716 13410
rect 1650 13392 1666 13394
rect 193 13362 219 13392
rect 1619 13362 1666 13392
rect 122 13298 188 13314
rect 122 13264 138 13298
rect 172 13296 188 13298
rect 1650 13360 1666 13362
rect 1700 13360 1716 13394
rect 1650 13344 1716 13360
rect 172 13266 219 13296
rect 1619 13266 1645 13296
rect 172 13264 188 13266
rect 122 13248 188 13264
rect 1650 13202 1716 13218
rect 1650 13200 1666 13202
rect 193 13170 219 13200
rect 1619 13170 1666 13200
rect 122 13106 188 13122
rect 122 13072 138 13106
rect 172 13104 188 13106
rect 1650 13168 1666 13170
rect 1700 13168 1716 13202
rect 1650 13152 1716 13168
rect 172 13074 219 13104
rect 1619 13074 1645 13104
rect 172 13072 188 13074
rect 122 13056 188 13072
rect 1650 13010 1716 13026
rect 1650 13008 1666 13010
rect 193 12978 219 13008
rect 1619 12978 1666 13008
rect 122 12914 188 12930
rect 122 12880 138 12914
rect 172 12912 188 12914
rect 1650 12976 1666 12978
rect 1700 12976 1716 13010
rect 1650 12960 1716 12976
rect 172 12882 219 12912
rect 1619 12882 1645 12912
rect 172 12880 188 12882
rect 122 12864 188 12880
rect 1650 12818 1716 12834
rect 1650 12816 1666 12818
rect 193 12786 219 12816
rect 1619 12786 1666 12816
rect 122 12722 188 12738
rect 122 12688 138 12722
rect 172 12720 188 12722
rect 1650 12784 1666 12786
rect 1700 12784 1716 12818
rect 1650 12768 1716 12784
rect 172 12690 219 12720
rect 1619 12690 1645 12720
rect 172 12688 188 12690
rect 122 12672 188 12688
rect 1650 12626 1716 12642
rect 1650 12624 1666 12626
rect 193 12594 219 12624
rect 1619 12594 1666 12624
rect 122 12530 188 12546
rect 122 12496 138 12530
rect 172 12528 188 12530
rect 1650 12592 1666 12594
rect 1700 12592 1716 12626
rect 1650 12576 1716 12592
rect 172 12498 219 12528
rect 1619 12498 1645 12528
rect 172 12496 188 12498
rect 122 12480 188 12496
rect 1650 12434 1716 12450
rect 1650 12432 1666 12434
rect 193 12402 219 12432
rect 1619 12402 1666 12432
rect 122 12338 188 12354
rect 122 12304 138 12338
rect 172 12336 188 12338
rect 1650 12400 1666 12402
rect 1700 12400 1716 12434
rect 1650 12384 1716 12400
rect 172 12306 219 12336
rect 1619 12306 1645 12336
rect 172 12304 188 12306
rect 122 12288 188 12304
rect 1650 12242 1716 12258
rect 1650 12240 1666 12242
rect 193 12210 219 12240
rect 1619 12210 1666 12240
rect 122 12146 188 12162
rect 122 12112 138 12146
rect 172 12144 188 12146
rect 1650 12208 1666 12210
rect 1700 12208 1716 12242
rect 1650 12192 1716 12208
rect 172 12114 219 12144
rect 1619 12114 1645 12144
rect 172 12112 188 12114
rect 122 12096 188 12112
rect 1650 12050 1716 12066
rect 1650 12048 1666 12050
rect 193 12018 219 12048
rect 1619 12018 1666 12048
rect 122 11954 188 11970
rect 122 11920 138 11954
rect 172 11952 188 11954
rect 1650 12016 1666 12018
rect 1700 12016 1716 12050
rect 1650 12000 1716 12016
rect 172 11922 219 11952
rect 1619 11922 1645 11952
rect 172 11920 188 11922
rect 122 11904 188 11920
rect 1650 11858 1716 11874
rect 1650 11856 1666 11858
rect 193 11826 219 11856
rect 1619 11826 1666 11856
rect 122 11762 188 11778
rect 122 11728 138 11762
rect 172 11760 188 11762
rect 1650 11824 1666 11826
rect 1700 11824 1716 11858
rect 1650 11808 1716 11824
rect 172 11730 219 11760
rect 1619 11730 1645 11760
rect 172 11728 188 11730
rect 122 11712 188 11728
rect 1650 11666 1716 11682
rect 1650 11664 1666 11666
rect 193 11634 219 11664
rect 1619 11634 1666 11664
rect 122 11570 188 11586
rect 122 11536 138 11570
rect 172 11568 188 11570
rect 1650 11632 1666 11634
rect 1700 11632 1716 11666
rect 1650 11616 1716 11632
rect 172 11538 219 11568
rect 1619 11538 1645 11568
rect 172 11536 188 11538
rect 122 11520 188 11536
rect 1650 11474 1716 11490
rect 1650 11472 1666 11474
rect 193 11442 219 11472
rect 1619 11442 1666 11472
rect 122 11378 188 11394
rect 122 11344 138 11378
rect 172 11376 188 11378
rect 1650 11440 1666 11442
rect 1700 11440 1716 11474
rect 1650 11424 1716 11440
rect 172 11346 219 11376
rect 1619 11346 1645 11376
rect 172 11344 188 11346
rect 122 11328 188 11344
rect 1650 11282 1716 11298
rect 1650 11280 1666 11282
rect 193 11250 219 11280
rect 1619 11250 1666 11280
rect 122 11186 188 11202
rect 122 11152 138 11186
rect 172 11184 188 11186
rect 1650 11248 1666 11250
rect 1700 11248 1716 11282
rect 1650 11232 1716 11248
rect 172 11154 219 11184
rect 1619 11154 1645 11184
rect 172 11152 188 11154
rect 122 11136 188 11152
rect 1650 11090 1716 11106
rect 1650 11088 1666 11090
rect 193 11058 219 11088
rect 1619 11058 1666 11088
rect 122 10994 188 11010
rect 122 10960 138 10994
rect 172 10992 188 10994
rect 1650 11056 1666 11058
rect 1700 11056 1716 11090
rect 1650 11040 1716 11056
rect 172 10962 219 10992
rect 1619 10962 1645 10992
rect 172 10960 188 10962
rect 122 10944 188 10960
rect 1650 10898 1716 10914
rect 1650 10896 1666 10898
rect 193 10866 219 10896
rect 1619 10866 1666 10896
rect 122 10802 188 10818
rect 122 10768 138 10802
rect 172 10800 188 10802
rect 1650 10864 1666 10866
rect 1700 10864 1716 10898
rect 1650 10848 1716 10864
rect 172 10770 219 10800
rect 1619 10770 1645 10800
rect 172 10768 188 10770
rect 122 10752 188 10768
rect 1650 10706 1716 10722
rect 1650 10704 1666 10706
rect 193 10674 219 10704
rect 1619 10674 1666 10704
rect 122 10610 188 10626
rect 122 10576 138 10610
rect 172 10608 188 10610
rect 1650 10672 1666 10674
rect 1700 10672 1716 10706
rect 1650 10656 1716 10672
rect 172 10578 219 10608
rect 1619 10578 1645 10608
rect 172 10576 188 10578
rect 122 10560 188 10576
rect 1650 10514 1716 10530
rect 1650 10512 1666 10514
rect 193 10482 219 10512
rect 1619 10482 1666 10512
rect 122 10418 188 10434
rect 122 10384 138 10418
rect 172 10416 188 10418
rect 1650 10480 1666 10482
rect 1700 10480 1716 10514
rect 1650 10464 1716 10480
rect 172 10386 219 10416
rect 1619 10386 1645 10416
rect 172 10384 188 10386
rect 122 10368 188 10384
rect 1650 10322 1716 10338
rect 1650 10320 1666 10322
rect 193 10290 219 10320
rect 1619 10290 1666 10320
rect 122 10226 188 10242
rect 122 10192 138 10226
rect 172 10224 188 10226
rect 1650 10288 1666 10290
rect 1700 10288 1716 10322
rect 1650 10272 1716 10288
rect 172 10194 219 10224
rect 1619 10194 1645 10224
rect 172 10192 188 10194
rect 122 10176 188 10192
rect 1650 10130 1716 10146
rect 1650 10128 1666 10130
rect 193 10098 219 10128
rect 1619 10098 1666 10128
rect 122 10034 188 10050
rect 122 10000 138 10034
rect 172 10032 188 10034
rect 1650 10096 1666 10098
rect 1700 10096 1716 10130
rect 1650 10080 1716 10096
rect 172 10002 219 10032
rect 1619 10002 1645 10032
rect 172 10000 188 10002
rect 122 9984 188 10000
rect 1650 9938 1716 9954
rect 1650 9936 1666 9938
rect 193 9906 219 9936
rect 1619 9906 1666 9936
rect 122 9842 188 9858
rect 122 9808 138 9842
rect 172 9840 188 9842
rect 1650 9904 1666 9906
rect 1700 9904 1716 9938
rect 1650 9888 1716 9904
rect 172 9810 219 9840
rect 1619 9810 1645 9840
rect 172 9808 188 9810
rect 122 9792 188 9808
rect 1650 9746 1716 9762
rect 1650 9744 1666 9746
rect 193 9714 219 9744
rect 1619 9714 1666 9744
rect 122 9650 188 9666
rect 122 9616 138 9650
rect 172 9648 188 9650
rect 1650 9712 1666 9714
rect 1700 9712 1716 9746
rect 1650 9696 1716 9712
rect 172 9618 219 9648
rect 1619 9618 1645 9648
rect 172 9616 188 9618
rect 122 9600 188 9616
rect 1650 9554 1716 9570
rect 1650 9552 1666 9554
rect 193 9522 219 9552
rect 1619 9522 1666 9552
rect 122 9458 188 9474
rect 122 9424 138 9458
rect 172 9456 188 9458
rect 1650 9520 1666 9522
rect 1700 9520 1716 9554
rect 1650 9504 1716 9520
rect 172 9426 219 9456
rect 1619 9426 1645 9456
rect 172 9424 188 9426
rect 122 9408 188 9424
rect 1650 9362 1716 9378
rect 1650 9360 1666 9362
rect 193 9330 219 9360
rect 1619 9330 1666 9360
rect 122 9266 188 9282
rect 122 9232 138 9266
rect 172 9264 188 9266
rect 1650 9328 1666 9330
rect 1700 9328 1716 9362
rect 1650 9312 1716 9328
rect 172 9234 219 9264
rect 1619 9234 1645 9264
rect 172 9232 188 9234
rect 122 9216 188 9232
rect 1650 9170 1716 9186
rect 1650 9168 1666 9170
rect 193 9138 219 9168
rect 1619 9138 1666 9168
rect 122 9074 188 9090
rect 122 9040 138 9074
rect 172 9072 188 9074
rect 1650 9136 1666 9138
rect 1700 9136 1716 9170
rect 1650 9120 1716 9136
rect 172 9042 219 9072
rect 1619 9042 1645 9072
rect 172 9040 188 9042
rect 122 9024 188 9040
rect 1650 8978 1716 8994
rect 1650 8976 1666 8978
rect 193 8946 219 8976
rect 1619 8946 1666 8976
rect 122 8882 188 8898
rect 122 8848 138 8882
rect 172 8880 188 8882
rect 1650 8944 1666 8946
rect 1700 8944 1716 8978
rect 1650 8928 1716 8944
rect 172 8850 219 8880
rect 1619 8850 1645 8880
rect 172 8848 188 8850
rect 122 8832 188 8848
rect 1650 8786 1716 8802
rect 1650 8784 1666 8786
rect 193 8754 219 8784
rect 1619 8754 1666 8784
rect 122 8690 188 8706
rect 122 8656 138 8690
rect 172 8688 188 8690
rect 1650 8752 1666 8754
rect 1700 8752 1716 8786
rect 1650 8736 1716 8752
rect 172 8658 219 8688
rect 1619 8658 1645 8688
rect 172 8656 188 8658
rect 122 8640 188 8656
rect 1650 8594 1716 8610
rect 1650 8592 1666 8594
rect 193 8562 219 8592
rect 1619 8562 1666 8592
rect 122 8498 188 8514
rect 122 8464 138 8498
rect 172 8496 188 8498
rect 1650 8560 1666 8562
rect 1700 8560 1716 8594
rect 1650 8544 1716 8560
rect 172 8466 219 8496
rect 1619 8466 1645 8496
rect 172 8464 188 8466
rect 122 8448 188 8464
rect 1650 8402 1716 8418
rect 1650 8400 1666 8402
rect 193 8370 219 8400
rect 1619 8370 1666 8400
rect 122 8306 188 8322
rect 122 8272 138 8306
rect 172 8304 188 8306
rect 1650 8368 1666 8370
rect 1700 8368 1716 8402
rect 1650 8352 1716 8368
rect 172 8274 219 8304
rect 1619 8274 1645 8304
rect 172 8272 188 8274
rect 122 8256 188 8272
rect 1650 8210 1716 8226
rect 1650 8208 1666 8210
rect 193 8178 219 8208
rect 1619 8178 1666 8208
rect 122 8114 188 8130
rect 122 8080 138 8114
rect 172 8112 188 8114
rect 1650 8176 1666 8178
rect 1700 8176 1716 8210
rect 1650 8160 1716 8176
rect 172 8082 219 8112
rect 1619 8082 1645 8112
rect 172 8080 188 8082
rect 122 8064 188 8080
rect 1650 8018 1716 8034
rect 1650 8016 1666 8018
rect 193 7986 219 8016
rect 1619 7986 1666 8016
rect 122 7922 188 7938
rect 122 7888 138 7922
rect 172 7920 188 7922
rect 1650 7984 1666 7986
rect 1700 7984 1716 8018
rect 1650 7968 1716 7984
rect 172 7890 219 7920
rect 1619 7890 1645 7920
rect 172 7888 188 7890
rect 122 7872 188 7888
rect 1650 7826 1716 7842
rect 1650 7824 1666 7826
rect 193 7794 219 7824
rect 1619 7794 1666 7824
rect 122 7730 188 7746
rect 122 7696 138 7730
rect 172 7728 188 7730
rect 1650 7792 1666 7794
rect 1700 7792 1716 7826
rect 1650 7776 1716 7792
rect 172 7698 219 7728
rect 1619 7698 1645 7728
rect 172 7696 188 7698
rect 122 7680 188 7696
rect 1650 7634 1716 7650
rect 1650 7632 1666 7634
rect 193 7602 219 7632
rect 1619 7602 1666 7632
rect 122 7538 188 7554
rect 122 7504 138 7538
rect 172 7536 188 7538
rect 1650 7600 1666 7602
rect 1700 7600 1716 7634
rect 1650 7584 1716 7600
rect 172 7506 219 7536
rect 1619 7506 1645 7536
rect 172 7504 188 7506
rect 122 7488 188 7504
rect 1650 7442 1716 7458
rect 1650 7440 1666 7442
rect 193 7410 219 7440
rect 1619 7410 1666 7440
rect 122 7346 188 7362
rect 122 7312 138 7346
rect 172 7344 188 7346
rect 1650 7408 1666 7410
rect 1700 7408 1716 7442
rect 1650 7392 1716 7408
rect 172 7314 219 7344
rect 1619 7314 1645 7344
rect 172 7312 188 7314
rect 122 7296 188 7312
rect 1650 7250 1716 7266
rect 1650 7248 1666 7250
rect 193 7218 219 7248
rect 1619 7218 1666 7248
rect 122 7154 188 7170
rect 122 7120 138 7154
rect 172 7152 188 7154
rect 1650 7216 1666 7218
rect 1700 7216 1716 7250
rect 1650 7200 1716 7216
rect 172 7122 219 7152
rect 1619 7122 1645 7152
rect 172 7120 188 7122
rect 122 7104 188 7120
rect 1650 7058 1716 7074
rect 1650 7056 1666 7058
rect 193 7026 219 7056
rect 1619 7026 1666 7056
rect 122 6962 188 6978
rect 122 6928 138 6962
rect 172 6960 188 6962
rect 1650 7024 1666 7026
rect 1700 7024 1716 7058
rect 1650 7008 1716 7024
rect 172 6930 219 6960
rect 1619 6930 1645 6960
rect 172 6928 188 6930
rect 122 6912 188 6928
rect 1650 6866 1716 6882
rect 1650 6864 1666 6866
rect 193 6834 219 6864
rect 1619 6834 1666 6864
rect 122 6770 188 6786
rect 122 6736 138 6770
rect 172 6768 188 6770
rect 1650 6832 1666 6834
rect 1700 6832 1716 6866
rect 1650 6816 1716 6832
rect 172 6738 219 6768
rect 1619 6738 1645 6768
rect 172 6736 188 6738
rect 122 6720 188 6736
rect 1650 6674 1716 6690
rect 1650 6672 1666 6674
rect 193 6642 219 6672
rect 1619 6642 1666 6672
rect 122 6578 188 6594
rect 122 6544 138 6578
rect 172 6576 188 6578
rect 1650 6640 1666 6642
rect 1700 6640 1716 6674
rect 1650 6624 1716 6640
rect 172 6546 219 6576
rect 1619 6546 1645 6576
rect 172 6544 188 6546
rect 122 6528 188 6544
rect 1650 6482 1716 6498
rect 1650 6480 1666 6482
rect 193 6450 219 6480
rect 1619 6450 1666 6480
rect 122 6386 188 6402
rect 122 6352 138 6386
rect 172 6384 188 6386
rect 1650 6448 1666 6450
rect 1700 6448 1716 6482
rect 1650 6432 1716 6448
rect 172 6354 219 6384
rect 1619 6354 1645 6384
rect 172 6352 188 6354
rect 122 6336 188 6352
rect 1650 6290 1716 6306
rect 1650 6288 1666 6290
rect 193 6258 219 6288
rect 1619 6258 1666 6288
rect 122 6194 188 6210
rect 122 6160 138 6194
rect 172 6192 188 6194
rect 1650 6256 1666 6258
rect 1700 6256 1716 6290
rect 1650 6240 1716 6256
rect 172 6162 219 6192
rect 1619 6162 1645 6192
rect 172 6160 188 6162
rect 122 6144 188 6160
rect 1650 6098 1716 6114
rect 1650 6096 1666 6098
rect 193 6066 219 6096
rect 1619 6066 1666 6096
rect 122 6002 188 6018
rect 122 5968 138 6002
rect 172 6000 188 6002
rect 1650 6064 1666 6066
rect 1700 6064 1716 6098
rect 1650 6048 1716 6064
rect 172 5970 219 6000
rect 1619 5970 1645 6000
rect 172 5968 188 5970
rect 122 5952 188 5968
rect 1650 5906 1716 5922
rect 1650 5904 1666 5906
rect 193 5874 219 5904
rect 1619 5874 1666 5904
rect 122 5810 188 5826
rect 122 5776 138 5810
rect 172 5808 188 5810
rect 1650 5872 1666 5874
rect 1700 5872 1716 5906
rect 1650 5856 1716 5872
rect 172 5778 219 5808
rect 1619 5778 1645 5808
rect 172 5776 188 5778
rect 122 5760 188 5776
rect 1650 5714 1716 5730
rect 1650 5712 1666 5714
rect 193 5682 219 5712
rect 1619 5682 1666 5712
rect 122 5618 188 5634
rect 122 5584 138 5618
rect 172 5616 188 5618
rect 1650 5680 1666 5682
rect 1700 5680 1716 5714
rect 1650 5664 1716 5680
rect 172 5586 219 5616
rect 1619 5586 1645 5616
rect 172 5584 188 5586
rect 122 5568 188 5584
rect 1650 5522 1716 5538
rect 1650 5520 1666 5522
rect 193 5490 219 5520
rect 1619 5490 1666 5520
rect 122 5426 188 5442
rect 122 5392 138 5426
rect 172 5424 188 5426
rect 1650 5488 1666 5490
rect 1700 5488 1716 5522
rect 1650 5472 1716 5488
rect 172 5394 219 5424
rect 1619 5394 1645 5424
rect 172 5392 188 5394
rect 122 5376 188 5392
rect 1650 5330 1716 5346
rect 1650 5328 1666 5330
rect 193 5298 219 5328
rect 1619 5298 1666 5328
rect 122 5234 188 5250
rect 122 5200 138 5234
rect 172 5232 188 5234
rect 1650 5296 1666 5298
rect 1700 5296 1716 5330
rect 1650 5280 1716 5296
rect 172 5202 219 5232
rect 1619 5202 1645 5232
rect 172 5200 188 5202
rect 122 5184 188 5200
rect 1650 5138 1716 5154
rect 1650 5136 1666 5138
rect 193 5106 219 5136
rect 1619 5106 1666 5136
rect 122 5042 188 5058
rect 122 5008 138 5042
rect 172 5040 188 5042
rect 1650 5104 1666 5106
rect 1700 5104 1716 5138
rect 1650 5088 1716 5104
rect 172 5010 219 5040
rect 1619 5010 1645 5040
rect 172 5008 188 5010
rect 122 4992 188 5008
rect 1650 4946 1716 4962
rect 1650 4944 1666 4946
rect 193 4914 219 4944
rect 1619 4914 1666 4944
rect 122 4850 188 4866
rect 122 4816 138 4850
rect 172 4848 188 4850
rect 1650 4912 1666 4914
rect 1700 4912 1716 4946
rect 1650 4896 1716 4912
rect 172 4818 219 4848
rect 1619 4818 1645 4848
rect 172 4816 188 4818
rect 122 4800 188 4816
rect 1650 4754 1716 4770
rect 1650 4752 1666 4754
rect 193 4722 219 4752
rect 1619 4722 1666 4752
rect 122 4658 188 4674
rect 122 4624 138 4658
rect 172 4656 188 4658
rect 1650 4720 1666 4722
rect 1700 4720 1716 4754
rect 1650 4704 1716 4720
rect 172 4626 219 4656
rect 1619 4626 1645 4656
rect 172 4624 188 4626
rect 122 4608 188 4624
rect 1650 4562 1716 4578
rect 1650 4560 1666 4562
rect 193 4530 219 4560
rect 1619 4530 1666 4560
rect 122 4466 188 4482
rect 122 4432 138 4466
rect 172 4464 188 4466
rect 1650 4528 1666 4530
rect 1700 4528 1716 4562
rect 1650 4512 1716 4528
rect 172 4434 219 4464
rect 1619 4434 1645 4464
rect 172 4432 188 4434
rect 122 4416 188 4432
rect 1650 4370 1716 4386
rect 1650 4368 1666 4370
rect 193 4338 219 4368
rect 1619 4338 1666 4368
rect 122 4274 188 4290
rect 122 4240 138 4274
rect 172 4272 188 4274
rect 1650 4336 1666 4338
rect 1700 4336 1716 4370
rect 1650 4320 1716 4336
rect 172 4242 219 4272
rect 1619 4242 1645 4272
rect 172 4240 188 4242
rect 122 4224 188 4240
rect 1650 4178 1716 4194
rect 1650 4176 1666 4178
rect 193 4146 219 4176
rect 1619 4146 1666 4176
rect 122 4082 188 4098
rect 122 4048 138 4082
rect 172 4080 188 4082
rect 1650 4144 1666 4146
rect 1700 4144 1716 4178
rect 1650 4128 1716 4144
rect 172 4050 219 4080
rect 1619 4050 1645 4080
rect 172 4048 188 4050
rect 122 4032 188 4048
rect 1650 3986 1716 4002
rect 1650 3984 1666 3986
rect 193 3954 219 3984
rect 1619 3954 1666 3984
rect 122 3890 188 3906
rect 122 3856 138 3890
rect 172 3888 188 3890
rect 1650 3952 1666 3954
rect 1700 3952 1716 3986
rect 1650 3936 1716 3952
rect 172 3858 219 3888
rect 1619 3858 1645 3888
rect 172 3856 188 3858
rect 122 3840 188 3856
rect 1650 3794 1716 3810
rect 1650 3792 1666 3794
rect 193 3762 219 3792
rect 1619 3762 1666 3792
rect 122 3698 188 3714
rect 122 3664 138 3698
rect 172 3696 188 3698
rect 1650 3760 1666 3762
rect 1700 3760 1716 3794
rect 1650 3744 1716 3760
rect 172 3666 219 3696
rect 1619 3666 1645 3696
rect 172 3664 188 3666
rect 122 3648 188 3664
rect 1650 3602 1716 3618
rect 1650 3600 1666 3602
rect 193 3570 219 3600
rect 1619 3570 1666 3600
rect 122 3506 188 3522
rect 122 3472 138 3506
rect 172 3504 188 3506
rect 1650 3568 1666 3570
rect 1700 3568 1716 3602
rect 1650 3552 1716 3568
rect 172 3474 219 3504
rect 1619 3474 1645 3504
rect 172 3472 188 3474
rect 122 3456 188 3472
rect 1650 3410 1716 3426
rect 1650 3408 1666 3410
rect 193 3378 219 3408
rect 1619 3378 1666 3408
rect 122 3314 188 3330
rect 122 3280 138 3314
rect 172 3312 188 3314
rect 1650 3376 1666 3378
rect 1700 3376 1716 3410
rect 1650 3360 1716 3376
rect 172 3282 219 3312
rect 1619 3282 1645 3312
rect 172 3280 188 3282
rect 122 3264 188 3280
rect 1650 3218 1716 3234
rect 1650 3216 1666 3218
rect 193 3186 219 3216
rect 1619 3186 1666 3216
rect 122 3122 188 3138
rect 122 3088 138 3122
rect 172 3120 188 3122
rect 1650 3184 1666 3186
rect 1700 3184 1716 3218
rect 1650 3168 1716 3184
rect 172 3090 219 3120
rect 1619 3090 1645 3120
rect 172 3088 188 3090
rect 122 3072 188 3088
rect 1650 3026 1716 3042
rect 1650 3024 1666 3026
rect 193 2994 219 3024
rect 1619 2994 1666 3024
rect 122 2930 188 2946
rect 122 2896 138 2930
rect 172 2928 188 2930
rect 1650 2992 1666 2994
rect 1700 2992 1716 3026
rect 1650 2976 1716 2992
rect 172 2898 219 2928
rect 1619 2898 1645 2928
rect 172 2896 188 2898
rect 122 2880 188 2896
rect 1650 2834 1716 2850
rect 1650 2832 1666 2834
rect 193 2802 219 2832
rect 1619 2802 1666 2832
rect 122 2738 188 2754
rect 122 2704 138 2738
rect 172 2736 188 2738
rect 1650 2800 1666 2802
rect 1700 2800 1716 2834
rect 1650 2784 1716 2800
rect 172 2706 219 2736
rect 1619 2706 1645 2736
rect 172 2704 188 2706
rect 122 2688 188 2704
rect 1650 2642 1716 2658
rect 1650 2640 1666 2642
rect 193 2610 219 2640
rect 1619 2610 1666 2640
rect 122 2546 188 2562
rect 122 2512 138 2546
rect 172 2544 188 2546
rect 1650 2608 1666 2610
rect 1700 2608 1716 2642
rect 1650 2592 1716 2608
rect 172 2514 219 2544
rect 1619 2514 1645 2544
rect 172 2512 188 2514
rect 122 2496 188 2512
rect 1650 2450 1716 2466
rect 1650 2448 1666 2450
rect 193 2418 219 2448
rect 1619 2418 1666 2448
rect 122 2354 188 2370
rect 122 2320 138 2354
rect 172 2352 188 2354
rect 1650 2416 1666 2418
rect 1700 2416 1716 2450
rect 1650 2400 1716 2416
rect 172 2322 219 2352
rect 1619 2322 1645 2352
rect 172 2320 188 2322
rect 122 2304 188 2320
rect 1650 2258 1716 2274
rect 1650 2256 1666 2258
rect 193 2226 219 2256
rect 1619 2226 1666 2256
rect 122 2162 188 2178
rect 122 2128 138 2162
rect 172 2160 188 2162
rect 1650 2224 1666 2226
rect 1700 2224 1716 2258
rect 1650 2208 1716 2224
rect 172 2130 219 2160
rect 1619 2130 1645 2160
rect 172 2128 188 2130
rect 122 2112 188 2128
rect 1650 2066 1716 2082
rect 1650 2064 1666 2066
rect 193 2034 219 2064
rect 1619 2034 1666 2064
rect 122 1970 188 1986
rect 122 1936 138 1970
rect 172 1968 188 1970
rect 1650 2032 1666 2034
rect 1700 2032 1716 2066
rect 1650 2016 1716 2032
rect 172 1938 219 1968
rect 1619 1938 1645 1968
rect 172 1936 188 1938
rect 122 1920 188 1936
rect 1650 1874 1716 1890
rect 1650 1872 1666 1874
rect 193 1842 219 1872
rect 1619 1842 1666 1872
rect 122 1778 188 1794
rect 122 1744 138 1778
rect 172 1776 188 1778
rect 1650 1840 1666 1842
rect 1700 1840 1716 1874
rect 1650 1824 1716 1840
rect 172 1746 219 1776
rect 1619 1746 1645 1776
rect 172 1744 188 1746
rect 122 1728 188 1744
rect 1650 1682 1716 1698
rect 1650 1680 1666 1682
rect 193 1650 219 1680
rect 1619 1650 1666 1680
rect 122 1586 188 1602
rect 122 1552 138 1586
rect 172 1584 188 1586
rect 1650 1648 1666 1650
rect 1700 1648 1716 1682
rect 1650 1632 1716 1648
rect 172 1554 219 1584
rect 1619 1554 1645 1584
rect 172 1552 188 1554
rect 122 1536 188 1552
rect 1650 1490 1716 1506
rect 1650 1488 1666 1490
rect 193 1458 219 1488
rect 1619 1458 1666 1488
rect 122 1394 188 1410
rect 122 1360 138 1394
rect 172 1392 188 1394
rect 1650 1456 1666 1458
rect 1700 1456 1716 1490
rect 1650 1440 1716 1456
rect 172 1362 219 1392
rect 1619 1362 1645 1392
rect 172 1360 188 1362
rect 122 1344 188 1360
rect 1650 1298 1716 1314
rect 1650 1296 1666 1298
rect 193 1266 219 1296
rect 1619 1266 1666 1296
rect 122 1202 188 1218
rect 122 1168 138 1202
rect 172 1200 188 1202
rect 1650 1264 1666 1266
rect 1700 1264 1716 1298
rect 1650 1248 1716 1264
rect 172 1170 219 1200
rect 1619 1170 1645 1200
rect 172 1168 188 1170
rect 122 1152 188 1168
rect 1650 1106 1716 1122
rect 1650 1104 1666 1106
rect 193 1074 219 1104
rect 1619 1074 1666 1104
rect 122 1010 188 1026
rect 122 976 138 1010
rect 172 1008 188 1010
rect 1650 1072 1666 1074
rect 1700 1072 1716 1106
rect 1650 1056 1716 1072
rect 172 978 219 1008
rect 1619 978 1645 1008
rect 172 976 188 978
rect 122 960 188 976
rect 1650 914 1716 930
rect 1650 912 1666 914
rect 193 882 219 912
rect 1619 882 1666 912
rect 122 818 188 834
rect 122 784 138 818
rect 172 816 188 818
rect 1650 880 1666 882
rect 1700 880 1716 914
rect 1650 864 1716 880
rect 172 786 219 816
rect 1619 786 1645 816
rect 172 784 188 786
rect 122 768 188 784
rect 1650 722 1716 738
rect 1650 720 1666 722
rect 193 690 219 720
rect 1619 690 1666 720
rect 1650 688 1666 690
rect 1700 688 1716 722
rect 1650 672 1716 688
<< polycont >>
rect 138 21712 172 21746
rect 138 21520 172 21554
rect 1666 21616 1700 21650
rect 138 21328 172 21362
rect 1666 21424 1700 21458
rect 138 21136 172 21170
rect 1666 21232 1700 21266
rect 138 20944 172 20978
rect 1666 21040 1700 21074
rect 138 20752 172 20786
rect 1666 20848 1700 20882
rect 138 20560 172 20594
rect 1666 20656 1700 20690
rect 138 20368 172 20402
rect 1666 20464 1700 20498
rect 138 20176 172 20210
rect 1666 20272 1700 20306
rect 138 19984 172 20018
rect 1666 20080 1700 20114
rect 138 19792 172 19826
rect 1666 19888 1700 19922
rect 138 19600 172 19634
rect 1666 19696 1700 19730
rect 138 19408 172 19442
rect 1666 19504 1700 19538
rect 138 19216 172 19250
rect 1666 19312 1700 19346
rect 138 19024 172 19058
rect 1666 19120 1700 19154
rect 138 18832 172 18866
rect 1666 18928 1700 18962
rect 138 18640 172 18674
rect 1666 18736 1700 18770
rect 138 18448 172 18482
rect 1666 18544 1700 18578
rect 138 18256 172 18290
rect 1666 18352 1700 18386
rect 138 18064 172 18098
rect 1666 18160 1700 18194
rect 138 17872 172 17906
rect 1666 17968 1700 18002
rect 138 17680 172 17714
rect 1666 17776 1700 17810
rect 138 17488 172 17522
rect 1666 17584 1700 17618
rect 138 17296 172 17330
rect 1666 17392 1700 17426
rect 138 17104 172 17138
rect 1666 17200 1700 17234
rect 138 16912 172 16946
rect 1666 17008 1700 17042
rect 138 16720 172 16754
rect 1666 16816 1700 16850
rect 138 16528 172 16562
rect 1666 16624 1700 16658
rect 138 16336 172 16370
rect 1666 16432 1700 16466
rect 138 16144 172 16178
rect 1666 16240 1700 16274
rect 138 15952 172 15986
rect 1666 16048 1700 16082
rect 138 15760 172 15794
rect 1666 15856 1700 15890
rect 138 15568 172 15602
rect 1666 15664 1700 15698
rect 138 15376 172 15410
rect 1666 15472 1700 15506
rect 138 15184 172 15218
rect 1666 15280 1700 15314
rect 138 14992 172 15026
rect 1666 15088 1700 15122
rect 138 14800 172 14834
rect 1666 14896 1700 14930
rect 138 14608 172 14642
rect 1666 14704 1700 14738
rect 138 14416 172 14450
rect 1666 14512 1700 14546
rect 138 14224 172 14258
rect 1666 14320 1700 14354
rect 138 14032 172 14066
rect 1666 14128 1700 14162
rect 138 13840 172 13874
rect 1666 13936 1700 13970
rect 138 13648 172 13682
rect 1666 13744 1700 13778
rect 138 13456 172 13490
rect 1666 13552 1700 13586
rect 138 13264 172 13298
rect 1666 13360 1700 13394
rect 138 13072 172 13106
rect 1666 13168 1700 13202
rect 138 12880 172 12914
rect 1666 12976 1700 13010
rect 138 12688 172 12722
rect 1666 12784 1700 12818
rect 138 12496 172 12530
rect 1666 12592 1700 12626
rect 138 12304 172 12338
rect 1666 12400 1700 12434
rect 138 12112 172 12146
rect 1666 12208 1700 12242
rect 138 11920 172 11954
rect 1666 12016 1700 12050
rect 138 11728 172 11762
rect 1666 11824 1700 11858
rect 138 11536 172 11570
rect 1666 11632 1700 11666
rect 138 11344 172 11378
rect 1666 11440 1700 11474
rect 138 11152 172 11186
rect 1666 11248 1700 11282
rect 138 10960 172 10994
rect 1666 11056 1700 11090
rect 138 10768 172 10802
rect 1666 10864 1700 10898
rect 138 10576 172 10610
rect 1666 10672 1700 10706
rect 138 10384 172 10418
rect 1666 10480 1700 10514
rect 138 10192 172 10226
rect 1666 10288 1700 10322
rect 138 10000 172 10034
rect 1666 10096 1700 10130
rect 138 9808 172 9842
rect 1666 9904 1700 9938
rect 138 9616 172 9650
rect 1666 9712 1700 9746
rect 138 9424 172 9458
rect 1666 9520 1700 9554
rect 138 9232 172 9266
rect 1666 9328 1700 9362
rect 138 9040 172 9074
rect 1666 9136 1700 9170
rect 138 8848 172 8882
rect 1666 8944 1700 8978
rect 138 8656 172 8690
rect 1666 8752 1700 8786
rect 138 8464 172 8498
rect 1666 8560 1700 8594
rect 138 8272 172 8306
rect 1666 8368 1700 8402
rect 138 8080 172 8114
rect 1666 8176 1700 8210
rect 138 7888 172 7922
rect 1666 7984 1700 8018
rect 138 7696 172 7730
rect 1666 7792 1700 7826
rect 138 7504 172 7538
rect 1666 7600 1700 7634
rect 138 7312 172 7346
rect 1666 7408 1700 7442
rect 138 7120 172 7154
rect 1666 7216 1700 7250
rect 138 6928 172 6962
rect 1666 7024 1700 7058
rect 138 6736 172 6770
rect 1666 6832 1700 6866
rect 138 6544 172 6578
rect 1666 6640 1700 6674
rect 138 6352 172 6386
rect 1666 6448 1700 6482
rect 138 6160 172 6194
rect 1666 6256 1700 6290
rect 138 5968 172 6002
rect 1666 6064 1700 6098
rect 138 5776 172 5810
rect 1666 5872 1700 5906
rect 138 5584 172 5618
rect 1666 5680 1700 5714
rect 138 5392 172 5426
rect 1666 5488 1700 5522
rect 138 5200 172 5234
rect 1666 5296 1700 5330
rect 138 5008 172 5042
rect 1666 5104 1700 5138
rect 138 4816 172 4850
rect 1666 4912 1700 4946
rect 138 4624 172 4658
rect 1666 4720 1700 4754
rect 138 4432 172 4466
rect 1666 4528 1700 4562
rect 138 4240 172 4274
rect 1666 4336 1700 4370
rect 138 4048 172 4082
rect 1666 4144 1700 4178
rect 138 3856 172 3890
rect 1666 3952 1700 3986
rect 138 3664 172 3698
rect 1666 3760 1700 3794
rect 138 3472 172 3506
rect 1666 3568 1700 3602
rect 138 3280 172 3314
rect 1666 3376 1700 3410
rect 138 3088 172 3122
rect 1666 3184 1700 3218
rect 138 2896 172 2930
rect 1666 2992 1700 3026
rect 138 2704 172 2738
rect 1666 2800 1700 2834
rect 138 2512 172 2546
rect 1666 2608 1700 2642
rect 138 2320 172 2354
rect 1666 2416 1700 2450
rect 138 2128 172 2162
rect 1666 2224 1700 2258
rect 138 1936 172 1970
rect 1666 2032 1700 2066
rect 138 1744 172 1778
rect 1666 1840 1700 1874
rect 138 1552 172 1586
rect 1666 1648 1700 1682
rect 138 1360 172 1394
rect 1666 1456 1700 1490
rect 138 1168 172 1202
rect 1666 1264 1700 1298
rect 138 976 172 1010
rect 1666 1072 1700 1106
rect 138 784 172 818
rect 1666 880 1700 914
rect 1666 688 1700 722
<< locali >>
rect 36 21874 132 21908
rect 1706 21874 1802 21908
rect 36 21812 70 21874
rect 1768 21812 1802 21874
rect 138 21746 172 21762
rect 215 21760 231 21794
rect 1607 21760 1623 21794
rect 138 21696 172 21712
rect 215 21664 231 21698
rect 1607 21664 1623 21698
rect 1666 21650 1700 21666
rect 138 21554 172 21570
rect 215 21568 231 21602
rect 1607 21568 1623 21602
rect 1666 21600 1700 21616
rect 138 21504 172 21520
rect 215 21472 231 21506
rect 1607 21472 1623 21506
rect 1666 21458 1700 21474
rect 138 21362 172 21378
rect 215 21376 231 21410
rect 1607 21376 1623 21410
rect 1666 21408 1700 21424
rect 138 21312 172 21328
rect 215 21280 231 21314
rect 1607 21280 1623 21314
rect 1666 21266 1700 21282
rect 138 21170 172 21186
rect 215 21184 231 21218
rect 1607 21184 1623 21218
rect 1666 21216 1700 21232
rect 138 21120 172 21136
rect 215 21088 231 21122
rect 1607 21088 1623 21122
rect 1666 21074 1700 21090
rect 138 20978 172 20994
rect 215 20992 231 21026
rect 1607 20992 1623 21026
rect 1666 21024 1700 21040
rect 138 20928 172 20944
rect 215 20896 231 20930
rect 1607 20896 1623 20930
rect 1666 20882 1700 20898
rect 138 20786 172 20802
rect 215 20800 231 20834
rect 1607 20800 1623 20834
rect 1666 20832 1700 20848
rect 138 20736 172 20752
rect 215 20704 231 20738
rect 1607 20704 1623 20738
rect 1666 20690 1700 20706
rect 138 20594 172 20610
rect 215 20608 231 20642
rect 1607 20608 1623 20642
rect 1666 20640 1700 20656
rect 138 20544 172 20560
rect 215 20512 231 20546
rect 1607 20512 1623 20546
rect 1666 20498 1700 20514
rect 138 20402 172 20418
rect 215 20416 231 20450
rect 1607 20416 1623 20450
rect 1666 20448 1700 20464
rect 138 20352 172 20368
rect 215 20320 231 20354
rect 1607 20320 1623 20354
rect 1666 20306 1700 20322
rect 138 20210 172 20226
rect 215 20224 231 20258
rect 1607 20224 1623 20258
rect 1666 20256 1700 20272
rect 138 20160 172 20176
rect 215 20128 231 20162
rect 1607 20128 1623 20162
rect 1666 20114 1700 20130
rect 138 20018 172 20034
rect 215 20032 231 20066
rect 1607 20032 1623 20066
rect 1666 20064 1700 20080
rect 138 19968 172 19984
rect 215 19936 231 19970
rect 1607 19936 1623 19970
rect 1666 19922 1700 19938
rect 138 19826 172 19842
rect 215 19840 231 19874
rect 1607 19840 1623 19874
rect 1666 19872 1700 19888
rect 138 19776 172 19792
rect 215 19744 231 19778
rect 1607 19744 1623 19778
rect 1666 19730 1700 19746
rect 138 19634 172 19650
rect 215 19648 231 19682
rect 1607 19648 1623 19682
rect 1666 19680 1700 19696
rect 138 19584 172 19600
rect 215 19552 231 19586
rect 1607 19552 1623 19586
rect 1666 19538 1700 19554
rect 138 19442 172 19458
rect 215 19456 231 19490
rect 1607 19456 1623 19490
rect 1666 19488 1700 19504
rect 138 19392 172 19408
rect 215 19360 231 19394
rect 1607 19360 1623 19394
rect 1666 19346 1700 19362
rect 138 19250 172 19266
rect 215 19264 231 19298
rect 1607 19264 1623 19298
rect 1666 19296 1700 19312
rect 138 19200 172 19216
rect 215 19168 231 19202
rect 1607 19168 1623 19202
rect 1666 19154 1700 19170
rect 138 19058 172 19074
rect 215 19072 231 19106
rect 1607 19072 1623 19106
rect 1666 19104 1700 19120
rect 138 19008 172 19024
rect 215 18976 231 19010
rect 1607 18976 1623 19010
rect 1666 18962 1700 18978
rect 138 18866 172 18882
rect 215 18880 231 18914
rect 1607 18880 1623 18914
rect 1666 18912 1700 18928
rect 138 18816 172 18832
rect 215 18784 231 18818
rect 1607 18784 1623 18818
rect 1666 18770 1700 18786
rect 138 18674 172 18690
rect 215 18688 231 18722
rect 1607 18688 1623 18722
rect 1666 18720 1700 18736
rect 138 18624 172 18640
rect 215 18592 231 18626
rect 1607 18592 1623 18626
rect 1666 18578 1700 18594
rect 138 18482 172 18498
rect 215 18496 231 18530
rect 1607 18496 1623 18530
rect 1666 18528 1700 18544
rect 138 18432 172 18448
rect 215 18400 231 18434
rect 1607 18400 1623 18434
rect 1666 18386 1700 18402
rect 138 18290 172 18306
rect 215 18304 231 18338
rect 1607 18304 1623 18338
rect 1666 18336 1700 18352
rect 138 18240 172 18256
rect 215 18208 231 18242
rect 1607 18208 1623 18242
rect 1666 18194 1700 18210
rect 138 18098 172 18114
rect 215 18112 231 18146
rect 1607 18112 1623 18146
rect 1666 18144 1700 18160
rect 138 18048 172 18064
rect 215 18016 231 18050
rect 1607 18016 1623 18050
rect 1666 18002 1700 18018
rect 138 17906 172 17922
rect 215 17920 231 17954
rect 1607 17920 1623 17954
rect 1666 17952 1700 17968
rect 138 17856 172 17872
rect 215 17824 231 17858
rect 1607 17824 1623 17858
rect 1666 17810 1700 17826
rect 138 17714 172 17730
rect 215 17728 231 17762
rect 1607 17728 1623 17762
rect 1666 17760 1700 17776
rect 138 17664 172 17680
rect 215 17632 231 17666
rect 1607 17632 1623 17666
rect 1666 17618 1700 17634
rect 138 17522 172 17538
rect 215 17536 231 17570
rect 1607 17536 1623 17570
rect 1666 17568 1700 17584
rect 138 17472 172 17488
rect 215 17440 231 17474
rect 1607 17440 1623 17474
rect 1666 17426 1700 17442
rect 138 17330 172 17346
rect 215 17344 231 17378
rect 1607 17344 1623 17378
rect 1666 17376 1700 17392
rect 138 17280 172 17296
rect 215 17248 231 17282
rect 1607 17248 1623 17282
rect 1666 17234 1700 17250
rect 138 17138 172 17154
rect 215 17152 231 17186
rect 1607 17152 1623 17186
rect 1666 17184 1700 17200
rect 138 17088 172 17104
rect 215 17056 231 17090
rect 1607 17056 1623 17090
rect 1666 17042 1700 17058
rect 138 16946 172 16962
rect 215 16960 231 16994
rect 1607 16960 1623 16994
rect 1666 16992 1700 17008
rect 138 16896 172 16912
rect 215 16864 231 16898
rect 1607 16864 1623 16898
rect 1666 16850 1700 16866
rect 138 16754 172 16770
rect 215 16768 231 16802
rect 1607 16768 1623 16802
rect 1666 16800 1700 16816
rect 138 16704 172 16720
rect 215 16672 231 16706
rect 1607 16672 1623 16706
rect 1666 16658 1700 16674
rect 138 16562 172 16578
rect 215 16576 231 16610
rect 1607 16576 1623 16610
rect 1666 16608 1700 16624
rect 138 16512 172 16528
rect 215 16480 231 16514
rect 1607 16480 1623 16514
rect 1666 16466 1700 16482
rect 138 16370 172 16386
rect 215 16384 231 16418
rect 1607 16384 1623 16418
rect 1666 16416 1700 16432
rect 138 16320 172 16336
rect 215 16288 231 16322
rect 1607 16288 1623 16322
rect 1666 16274 1700 16290
rect 138 16178 172 16194
rect 215 16192 231 16226
rect 1607 16192 1623 16226
rect 1666 16224 1700 16240
rect 138 16128 172 16144
rect 215 16096 231 16130
rect 1607 16096 1623 16130
rect 1666 16082 1700 16098
rect 138 15986 172 16002
rect 215 16000 231 16034
rect 1607 16000 1623 16034
rect 1666 16032 1700 16048
rect 138 15936 172 15952
rect 215 15904 231 15938
rect 1607 15904 1623 15938
rect 1666 15890 1700 15906
rect 138 15794 172 15810
rect 215 15808 231 15842
rect 1607 15808 1623 15842
rect 1666 15840 1700 15856
rect 138 15744 172 15760
rect 215 15712 231 15746
rect 1607 15712 1623 15746
rect 1666 15698 1700 15714
rect 138 15602 172 15618
rect 215 15616 231 15650
rect 1607 15616 1623 15650
rect 1666 15648 1700 15664
rect 138 15552 172 15568
rect 215 15520 231 15554
rect 1607 15520 1623 15554
rect 1666 15506 1700 15522
rect 138 15410 172 15426
rect 215 15424 231 15458
rect 1607 15424 1623 15458
rect 1666 15456 1700 15472
rect 138 15360 172 15376
rect 215 15328 231 15362
rect 1607 15328 1623 15362
rect 1666 15314 1700 15330
rect 138 15218 172 15234
rect 215 15232 231 15266
rect 1607 15232 1623 15266
rect 1666 15264 1700 15280
rect 138 15168 172 15184
rect 215 15136 231 15170
rect 1607 15136 1623 15170
rect 1666 15122 1700 15138
rect 138 15026 172 15042
rect 215 15040 231 15074
rect 1607 15040 1623 15074
rect 1666 15072 1700 15088
rect 138 14976 172 14992
rect 215 14944 231 14978
rect 1607 14944 1623 14978
rect 1666 14930 1700 14946
rect 138 14834 172 14850
rect 215 14848 231 14882
rect 1607 14848 1623 14882
rect 1666 14880 1700 14896
rect 138 14784 172 14800
rect 215 14752 231 14786
rect 1607 14752 1623 14786
rect 1666 14738 1700 14754
rect 138 14642 172 14658
rect 215 14656 231 14690
rect 1607 14656 1623 14690
rect 1666 14688 1700 14704
rect 138 14592 172 14608
rect 215 14560 231 14594
rect 1607 14560 1623 14594
rect 1666 14546 1700 14562
rect 138 14450 172 14466
rect 215 14464 231 14498
rect 1607 14464 1623 14498
rect 1666 14496 1700 14512
rect 138 14400 172 14416
rect 215 14368 231 14402
rect 1607 14368 1623 14402
rect 1666 14354 1700 14370
rect 138 14258 172 14274
rect 215 14272 231 14306
rect 1607 14272 1623 14306
rect 1666 14304 1700 14320
rect 138 14208 172 14224
rect 215 14176 231 14210
rect 1607 14176 1623 14210
rect 1666 14162 1700 14178
rect 138 14066 172 14082
rect 215 14080 231 14114
rect 1607 14080 1623 14114
rect 1666 14112 1700 14128
rect 138 14016 172 14032
rect 215 13984 231 14018
rect 1607 13984 1623 14018
rect 1666 13970 1700 13986
rect 138 13874 172 13890
rect 215 13888 231 13922
rect 1607 13888 1623 13922
rect 1666 13920 1700 13936
rect 138 13824 172 13840
rect 215 13792 231 13826
rect 1607 13792 1623 13826
rect 1666 13778 1700 13794
rect 138 13682 172 13698
rect 215 13696 231 13730
rect 1607 13696 1623 13730
rect 1666 13728 1700 13744
rect 138 13632 172 13648
rect 215 13600 231 13634
rect 1607 13600 1623 13634
rect 1666 13586 1700 13602
rect 138 13490 172 13506
rect 215 13504 231 13538
rect 1607 13504 1623 13538
rect 1666 13536 1700 13552
rect 138 13440 172 13456
rect 215 13408 231 13442
rect 1607 13408 1623 13442
rect 1666 13394 1700 13410
rect 138 13298 172 13314
rect 215 13312 231 13346
rect 1607 13312 1623 13346
rect 1666 13344 1700 13360
rect 138 13248 172 13264
rect 215 13216 231 13250
rect 1607 13216 1623 13250
rect 1666 13202 1700 13218
rect 138 13106 172 13122
rect 215 13120 231 13154
rect 1607 13120 1623 13154
rect 1666 13152 1700 13168
rect 138 13056 172 13072
rect 215 13024 231 13058
rect 1607 13024 1623 13058
rect 1666 13010 1700 13026
rect 138 12914 172 12930
rect 215 12928 231 12962
rect 1607 12928 1623 12962
rect 1666 12960 1700 12976
rect 138 12864 172 12880
rect 215 12832 231 12866
rect 1607 12832 1623 12866
rect 1666 12818 1700 12834
rect 138 12722 172 12738
rect 215 12736 231 12770
rect 1607 12736 1623 12770
rect 1666 12768 1700 12784
rect 138 12672 172 12688
rect 215 12640 231 12674
rect 1607 12640 1623 12674
rect 1666 12626 1700 12642
rect 138 12530 172 12546
rect 215 12544 231 12578
rect 1607 12544 1623 12578
rect 1666 12576 1700 12592
rect 138 12480 172 12496
rect 215 12448 231 12482
rect 1607 12448 1623 12482
rect 1666 12434 1700 12450
rect 138 12338 172 12354
rect 215 12352 231 12386
rect 1607 12352 1623 12386
rect 1666 12384 1700 12400
rect 138 12288 172 12304
rect 215 12256 231 12290
rect 1607 12256 1623 12290
rect 1666 12242 1700 12258
rect 138 12146 172 12162
rect 215 12160 231 12194
rect 1607 12160 1623 12194
rect 1666 12192 1700 12208
rect 138 12096 172 12112
rect 215 12064 231 12098
rect 1607 12064 1623 12098
rect 1666 12050 1700 12066
rect 138 11954 172 11970
rect 215 11968 231 12002
rect 1607 11968 1623 12002
rect 1666 12000 1700 12016
rect 138 11904 172 11920
rect 215 11872 231 11906
rect 1607 11872 1623 11906
rect 1666 11858 1700 11874
rect 138 11762 172 11778
rect 215 11776 231 11810
rect 1607 11776 1623 11810
rect 1666 11808 1700 11824
rect 138 11712 172 11728
rect 215 11680 231 11714
rect 1607 11680 1623 11714
rect 1666 11666 1700 11682
rect 138 11570 172 11586
rect 215 11584 231 11618
rect 1607 11584 1623 11618
rect 1666 11616 1700 11632
rect 138 11520 172 11536
rect 215 11488 231 11522
rect 1607 11488 1623 11522
rect 1666 11474 1700 11490
rect 138 11378 172 11394
rect 215 11392 231 11426
rect 1607 11392 1623 11426
rect 1666 11424 1700 11440
rect 138 11328 172 11344
rect 215 11296 231 11330
rect 1607 11296 1623 11330
rect 1666 11282 1700 11298
rect 138 11186 172 11202
rect 215 11200 231 11234
rect 1607 11200 1623 11234
rect 1666 11232 1700 11248
rect 138 11136 172 11152
rect 215 11104 231 11138
rect 1607 11104 1623 11138
rect 1666 11090 1700 11106
rect 138 10994 172 11010
rect 215 11008 231 11042
rect 1607 11008 1623 11042
rect 1666 11040 1700 11056
rect 138 10944 172 10960
rect 215 10912 231 10946
rect 1607 10912 1623 10946
rect 1666 10898 1700 10914
rect 138 10802 172 10818
rect 215 10816 231 10850
rect 1607 10816 1623 10850
rect 1666 10848 1700 10864
rect 138 10752 172 10768
rect 215 10720 231 10754
rect 1607 10720 1623 10754
rect 1666 10706 1700 10722
rect 138 10610 172 10626
rect 215 10624 231 10658
rect 1607 10624 1623 10658
rect 1666 10656 1700 10672
rect 138 10560 172 10576
rect 215 10528 231 10562
rect 1607 10528 1623 10562
rect 1666 10514 1700 10530
rect 138 10418 172 10434
rect 215 10432 231 10466
rect 1607 10432 1623 10466
rect 1666 10464 1700 10480
rect 138 10368 172 10384
rect 215 10336 231 10370
rect 1607 10336 1623 10370
rect 1666 10322 1700 10338
rect 138 10226 172 10242
rect 215 10240 231 10274
rect 1607 10240 1623 10274
rect 1666 10272 1700 10288
rect 138 10176 172 10192
rect 215 10144 231 10178
rect 1607 10144 1623 10178
rect 1666 10130 1700 10146
rect 138 10034 172 10050
rect 215 10048 231 10082
rect 1607 10048 1623 10082
rect 1666 10080 1700 10096
rect 138 9984 172 10000
rect 215 9952 231 9986
rect 1607 9952 1623 9986
rect 1666 9938 1700 9954
rect 138 9842 172 9858
rect 215 9856 231 9890
rect 1607 9856 1623 9890
rect 1666 9888 1700 9904
rect 138 9792 172 9808
rect 215 9760 231 9794
rect 1607 9760 1623 9794
rect 1666 9746 1700 9762
rect 138 9650 172 9666
rect 215 9664 231 9698
rect 1607 9664 1623 9698
rect 1666 9696 1700 9712
rect 138 9600 172 9616
rect 215 9568 231 9602
rect 1607 9568 1623 9602
rect 1666 9554 1700 9570
rect 138 9458 172 9474
rect 215 9472 231 9506
rect 1607 9472 1623 9506
rect 1666 9504 1700 9520
rect 138 9408 172 9424
rect 215 9376 231 9410
rect 1607 9376 1623 9410
rect 1666 9362 1700 9378
rect 138 9266 172 9282
rect 215 9280 231 9314
rect 1607 9280 1623 9314
rect 1666 9312 1700 9328
rect 138 9216 172 9232
rect 215 9184 231 9218
rect 1607 9184 1623 9218
rect 1666 9170 1700 9186
rect 138 9074 172 9090
rect 215 9088 231 9122
rect 1607 9088 1623 9122
rect 1666 9120 1700 9136
rect 138 9024 172 9040
rect 215 8992 231 9026
rect 1607 8992 1623 9026
rect 1666 8978 1700 8994
rect 138 8882 172 8898
rect 215 8896 231 8930
rect 1607 8896 1623 8930
rect 1666 8928 1700 8944
rect 138 8832 172 8848
rect 215 8800 231 8834
rect 1607 8800 1623 8834
rect 1666 8786 1700 8802
rect 138 8690 172 8706
rect 215 8704 231 8738
rect 1607 8704 1623 8738
rect 1666 8736 1700 8752
rect 138 8640 172 8656
rect 215 8608 231 8642
rect 1607 8608 1623 8642
rect 1666 8594 1700 8610
rect 138 8498 172 8514
rect 215 8512 231 8546
rect 1607 8512 1623 8546
rect 1666 8544 1700 8560
rect 138 8448 172 8464
rect 215 8416 231 8450
rect 1607 8416 1623 8450
rect 1666 8402 1700 8418
rect 138 8306 172 8322
rect 215 8320 231 8354
rect 1607 8320 1623 8354
rect 1666 8352 1700 8368
rect 138 8256 172 8272
rect 215 8224 231 8258
rect 1607 8224 1623 8258
rect 1666 8210 1700 8226
rect 138 8114 172 8130
rect 215 8128 231 8162
rect 1607 8128 1623 8162
rect 1666 8160 1700 8176
rect 138 8064 172 8080
rect 215 8032 231 8066
rect 1607 8032 1623 8066
rect 1666 8018 1700 8034
rect 138 7922 172 7938
rect 215 7936 231 7970
rect 1607 7936 1623 7970
rect 1666 7968 1700 7984
rect 138 7872 172 7888
rect 215 7840 231 7874
rect 1607 7840 1623 7874
rect 1666 7826 1700 7842
rect 138 7730 172 7746
rect 215 7744 231 7778
rect 1607 7744 1623 7778
rect 1666 7776 1700 7792
rect 138 7680 172 7696
rect 215 7648 231 7682
rect 1607 7648 1623 7682
rect 1666 7634 1700 7650
rect 138 7538 172 7554
rect 215 7552 231 7586
rect 1607 7552 1623 7586
rect 1666 7584 1700 7600
rect 138 7488 172 7504
rect 215 7456 231 7490
rect 1607 7456 1623 7490
rect 1666 7442 1700 7458
rect 138 7346 172 7362
rect 215 7360 231 7394
rect 1607 7360 1623 7394
rect 1666 7392 1700 7408
rect 138 7296 172 7312
rect 215 7264 231 7298
rect 1607 7264 1623 7298
rect 1666 7250 1700 7266
rect 138 7154 172 7170
rect 215 7168 231 7202
rect 1607 7168 1623 7202
rect 1666 7200 1700 7216
rect 138 7104 172 7120
rect 215 7072 231 7106
rect 1607 7072 1623 7106
rect 1666 7058 1700 7074
rect 138 6962 172 6978
rect 215 6976 231 7010
rect 1607 6976 1623 7010
rect 1666 7008 1700 7024
rect 138 6912 172 6928
rect 215 6880 231 6914
rect 1607 6880 1623 6914
rect 1666 6866 1700 6882
rect 138 6770 172 6786
rect 215 6784 231 6818
rect 1607 6784 1623 6818
rect 1666 6816 1700 6832
rect 138 6720 172 6736
rect 215 6688 231 6722
rect 1607 6688 1623 6722
rect 1666 6674 1700 6690
rect 138 6578 172 6594
rect 215 6592 231 6626
rect 1607 6592 1623 6626
rect 1666 6624 1700 6640
rect 138 6528 172 6544
rect 215 6496 231 6530
rect 1607 6496 1623 6530
rect 1666 6482 1700 6498
rect 138 6386 172 6402
rect 215 6400 231 6434
rect 1607 6400 1623 6434
rect 1666 6432 1700 6448
rect 138 6336 172 6352
rect 215 6304 231 6338
rect 1607 6304 1623 6338
rect 1666 6290 1700 6306
rect 138 6194 172 6210
rect 215 6208 231 6242
rect 1607 6208 1623 6242
rect 1666 6240 1700 6256
rect 138 6144 172 6160
rect 215 6112 231 6146
rect 1607 6112 1623 6146
rect 1666 6098 1700 6114
rect 138 6002 172 6018
rect 215 6016 231 6050
rect 1607 6016 1623 6050
rect 1666 6048 1700 6064
rect 138 5952 172 5968
rect 215 5920 231 5954
rect 1607 5920 1623 5954
rect 1666 5906 1700 5922
rect 138 5810 172 5826
rect 215 5824 231 5858
rect 1607 5824 1623 5858
rect 1666 5856 1700 5872
rect 138 5760 172 5776
rect 215 5728 231 5762
rect 1607 5728 1623 5762
rect 1666 5714 1700 5730
rect 138 5618 172 5634
rect 215 5632 231 5666
rect 1607 5632 1623 5666
rect 1666 5664 1700 5680
rect 138 5568 172 5584
rect 215 5536 231 5570
rect 1607 5536 1623 5570
rect 1666 5522 1700 5538
rect 138 5426 172 5442
rect 215 5440 231 5474
rect 1607 5440 1623 5474
rect 1666 5472 1700 5488
rect 138 5376 172 5392
rect 215 5344 231 5378
rect 1607 5344 1623 5378
rect 1666 5330 1700 5346
rect 138 5234 172 5250
rect 215 5248 231 5282
rect 1607 5248 1623 5282
rect 1666 5280 1700 5296
rect 138 5184 172 5200
rect 215 5152 231 5186
rect 1607 5152 1623 5186
rect 1666 5138 1700 5154
rect 138 5042 172 5058
rect 215 5056 231 5090
rect 1607 5056 1623 5090
rect 1666 5088 1700 5104
rect 138 4992 172 5008
rect 215 4960 231 4994
rect 1607 4960 1623 4994
rect 1666 4946 1700 4962
rect 138 4850 172 4866
rect 215 4864 231 4898
rect 1607 4864 1623 4898
rect 1666 4896 1700 4912
rect 138 4800 172 4816
rect 215 4768 231 4802
rect 1607 4768 1623 4802
rect 1666 4754 1700 4770
rect 138 4658 172 4674
rect 215 4672 231 4706
rect 1607 4672 1623 4706
rect 1666 4704 1700 4720
rect 138 4608 172 4624
rect 215 4576 231 4610
rect 1607 4576 1623 4610
rect 1666 4562 1700 4578
rect 138 4466 172 4482
rect 215 4480 231 4514
rect 1607 4480 1623 4514
rect 1666 4512 1700 4528
rect 138 4416 172 4432
rect 215 4384 231 4418
rect 1607 4384 1623 4418
rect 1666 4370 1700 4386
rect 138 4274 172 4290
rect 215 4288 231 4322
rect 1607 4288 1623 4322
rect 1666 4320 1700 4336
rect 138 4224 172 4240
rect 215 4192 231 4226
rect 1607 4192 1623 4226
rect 1666 4178 1700 4194
rect 138 4082 172 4098
rect 215 4096 231 4130
rect 1607 4096 1623 4130
rect 1666 4128 1700 4144
rect 138 4032 172 4048
rect 215 4000 231 4034
rect 1607 4000 1623 4034
rect 1666 3986 1700 4002
rect 138 3890 172 3906
rect 215 3904 231 3938
rect 1607 3904 1623 3938
rect 1666 3936 1700 3952
rect 138 3840 172 3856
rect 215 3808 231 3842
rect 1607 3808 1623 3842
rect 1666 3794 1700 3810
rect 138 3698 172 3714
rect 215 3712 231 3746
rect 1607 3712 1623 3746
rect 1666 3744 1700 3760
rect 138 3648 172 3664
rect 215 3616 231 3650
rect 1607 3616 1623 3650
rect 1666 3602 1700 3618
rect 138 3506 172 3522
rect 215 3520 231 3554
rect 1607 3520 1623 3554
rect 1666 3552 1700 3568
rect 138 3456 172 3472
rect 215 3424 231 3458
rect 1607 3424 1623 3458
rect 1666 3410 1700 3426
rect 138 3314 172 3330
rect 215 3328 231 3362
rect 1607 3328 1623 3362
rect 1666 3360 1700 3376
rect 138 3264 172 3280
rect 215 3232 231 3266
rect 1607 3232 1623 3266
rect 1666 3218 1700 3234
rect 138 3122 172 3138
rect 215 3136 231 3170
rect 1607 3136 1623 3170
rect 1666 3168 1700 3184
rect 138 3072 172 3088
rect 215 3040 231 3074
rect 1607 3040 1623 3074
rect 1666 3026 1700 3042
rect 138 2930 172 2946
rect 215 2944 231 2978
rect 1607 2944 1623 2978
rect 1666 2976 1700 2992
rect 138 2880 172 2896
rect 215 2848 231 2882
rect 1607 2848 1623 2882
rect 1666 2834 1700 2850
rect 138 2738 172 2754
rect 215 2752 231 2786
rect 1607 2752 1623 2786
rect 1666 2784 1700 2800
rect 138 2688 172 2704
rect 215 2656 231 2690
rect 1607 2656 1623 2690
rect 1666 2642 1700 2658
rect 138 2546 172 2562
rect 215 2560 231 2594
rect 1607 2560 1623 2594
rect 1666 2592 1700 2608
rect 138 2496 172 2512
rect 215 2464 231 2498
rect 1607 2464 1623 2498
rect 1666 2450 1700 2466
rect 138 2354 172 2370
rect 215 2368 231 2402
rect 1607 2368 1623 2402
rect 1666 2400 1700 2416
rect 138 2304 172 2320
rect 215 2272 231 2306
rect 1607 2272 1623 2306
rect 1666 2258 1700 2274
rect 138 2162 172 2178
rect 215 2176 231 2210
rect 1607 2176 1623 2210
rect 1666 2208 1700 2224
rect 138 2112 172 2128
rect 215 2080 231 2114
rect 1607 2080 1623 2114
rect 1666 2066 1700 2082
rect 138 1970 172 1986
rect 215 1984 231 2018
rect 1607 1984 1623 2018
rect 1666 2016 1700 2032
rect 138 1920 172 1936
rect 215 1888 231 1922
rect 1607 1888 1623 1922
rect 1666 1874 1700 1890
rect 138 1778 172 1794
rect 215 1792 231 1826
rect 1607 1792 1623 1826
rect 1666 1824 1700 1840
rect 138 1728 172 1744
rect 215 1696 231 1730
rect 1607 1696 1623 1730
rect 1666 1682 1700 1698
rect 138 1586 172 1602
rect 215 1600 231 1634
rect 1607 1600 1623 1634
rect 1666 1632 1700 1648
rect 138 1536 172 1552
rect 215 1504 231 1538
rect 1607 1504 1623 1538
rect 1666 1490 1700 1506
rect 138 1394 172 1410
rect 215 1408 231 1442
rect 1607 1408 1623 1442
rect 1666 1440 1700 1456
rect 138 1344 172 1360
rect 215 1312 231 1346
rect 1607 1312 1623 1346
rect 1666 1298 1700 1314
rect 138 1202 172 1218
rect 215 1216 231 1250
rect 1607 1216 1623 1250
rect 1666 1248 1700 1264
rect 138 1152 172 1168
rect 215 1120 231 1154
rect 1607 1120 1623 1154
rect 1666 1106 1700 1122
rect 138 1010 172 1026
rect 215 1024 231 1058
rect 1607 1024 1623 1058
rect 1666 1056 1700 1072
rect 138 960 172 976
rect 215 928 231 962
rect 1607 928 1623 962
rect 1666 914 1700 930
rect 138 818 172 834
rect 215 832 231 866
rect 1607 832 1623 866
rect 1666 864 1700 880
rect 138 768 172 784
rect 215 736 231 770
rect 1607 736 1623 770
rect 1666 722 1700 738
rect 215 640 231 674
rect 1607 640 1623 674
rect 1666 672 1700 688
rect 36 560 70 622
rect 1768 560 1802 622
rect 36 526 132 560
rect 1706 526 1802 560
<< viali >>
rect 328 21908 882 21932
rect 328 21874 882 21908
rect 328 21868 882 21874
rect 231 21760 1607 21794
rect 138 21712 172 21746
rect 231 21664 1607 21698
rect 1666 21616 1700 21650
rect 231 21568 1607 21602
rect 138 21520 172 21554
rect 231 21472 1607 21506
rect 1666 21424 1700 21458
rect 231 21376 1607 21410
rect 138 21328 172 21362
rect 231 21280 1607 21314
rect 1666 21232 1700 21266
rect 231 21184 1607 21218
rect 138 21136 172 21170
rect 231 21088 1607 21122
rect 1666 21040 1700 21074
rect 231 20992 1607 21026
rect 138 20944 172 20978
rect 231 20896 1607 20930
rect 1666 20848 1700 20882
rect 231 20800 1607 20834
rect 138 20752 172 20786
rect 231 20704 1607 20738
rect 1666 20656 1700 20690
rect 231 20608 1607 20642
rect 138 20560 172 20594
rect 231 20512 1607 20546
rect 1666 20464 1700 20498
rect 231 20416 1607 20450
rect 138 20368 172 20402
rect 231 20320 1607 20354
rect 1666 20272 1700 20306
rect 231 20224 1607 20258
rect 138 20176 172 20210
rect 231 20128 1607 20162
rect 1666 20080 1700 20114
rect 231 20032 1607 20066
rect 138 19984 172 20018
rect 231 19936 1607 19970
rect 1666 19888 1700 19922
rect 231 19840 1607 19874
rect 138 19792 172 19826
rect 231 19744 1607 19778
rect 1666 19696 1700 19730
rect 231 19648 1607 19682
rect 138 19600 172 19634
rect 231 19552 1607 19586
rect 1666 19504 1700 19538
rect 231 19456 1607 19490
rect 138 19408 172 19442
rect 231 19360 1607 19394
rect 1666 19312 1700 19346
rect 231 19264 1607 19298
rect 138 19216 172 19250
rect 231 19168 1607 19202
rect 1666 19120 1700 19154
rect 231 19072 1607 19106
rect 138 19024 172 19058
rect 231 18976 1607 19010
rect 1666 18928 1700 18962
rect 231 18880 1607 18914
rect 138 18832 172 18866
rect 231 18784 1607 18818
rect 1666 18736 1700 18770
rect 231 18688 1607 18722
rect 138 18640 172 18674
rect 231 18592 1607 18626
rect 1666 18544 1700 18578
rect 231 18496 1607 18530
rect 138 18448 172 18482
rect 231 18400 1607 18434
rect 1666 18352 1700 18386
rect 231 18304 1607 18338
rect 138 18256 172 18290
rect 231 18208 1607 18242
rect 1666 18160 1700 18194
rect 231 18112 1607 18146
rect 138 18064 172 18098
rect 231 18016 1607 18050
rect 1666 17968 1700 18002
rect 231 17920 1607 17954
rect 138 17872 172 17906
rect 231 17824 1607 17858
rect 1666 17776 1700 17810
rect 231 17728 1607 17762
rect 138 17680 172 17714
rect 231 17632 1607 17666
rect 1666 17584 1700 17618
rect 231 17536 1607 17570
rect 138 17488 172 17522
rect 231 17440 1607 17474
rect 1666 17392 1700 17426
rect 231 17344 1607 17378
rect 138 17296 172 17330
rect 231 17248 1607 17282
rect 1666 17200 1700 17234
rect 231 17152 1607 17186
rect 138 17104 172 17138
rect 231 17056 1607 17090
rect 1666 17008 1700 17042
rect 231 16960 1607 16994
rect 138 16912 172 16946
rect 231 16864 1607 16898
rect 1666 16816 1700 16850
rect 231 16768 1607 16802
rect 138 16720 172 16754
rect 231 16672 1607 16706
rect 1666 16624 1700 16658
rect 231 16576 1607 16610
rect 138 16528 172 16562
rect 231 16480 1607 16514
rect 1666 16432 1700 16466
rect 231 16384 1607 16418
rect 138 16336 172 16370
rect 231 16288 1607 16322
rect 1666 16240 1700 16274
rect 231 16192 1607 16226
rect 138 16144 172 16178
rect 231 16096 1607 16130
rect 1666 16048 1700 16082
rect 231 16000 1607 16034
rect 138 15952 172 15986
rect 231 15904 1607 15938
rect 1666 15856 1700 15890
rect 231 15808 1607 15842
rect 138 15760 172 15794
rect 231 15712 1607 15746
rect 1666 15664 1700 15698
rect 231 15616 1607 15650
rect 138 15568 172 15602
rect 231 15520 1607 15554
rect 1666 15472 1700 15506
rect 231 15424 1607 15458
rect 138 15376 172 15410
rect 231 15328 1607 15362
rect 1666 15280 1700 15314
rect 231 15232 1607 15266
rect 138 15184 172 15218
rect 231 15136 1607 15170
rect 1666 15088 1700 15122
rect 231 15040 1607 15074
rect 138 14992 172 15026
rect 231 14944 1607 14978
rect 1666 14896 1700 14930
rect 231 14848 1607 14882
rect 138 14800 172 14834
rect 231 14752 1607 14786
rect 1666 14704 1700 14738
rect 231 14656 1607 14690
rect 138 14608 172 14642
rect 231 14560 1607 14594
rect 1666 14512 1700 14546
rect 231 14464 1607 14498
rect 138 14416 172 14450
rect 231 14368 1607 14402
rect 1666 14320 1700 14354
rect 231 14272 1607 14306
rect 138 14224 172 14258
rect 231 14176 1607 14210
rect 1666 14128 1700 14162
rect 231 14080 1607 14114
rect 138 14032 172 14066
rect 231 13984 1607 14018
rect 1666 13936 1700 13970
rect 231 13888 1607 13922
rect 138 13840 172 13874
rect 231 13792 1607 13826
rect 1666 13744 1700 13778
rect 231 13696 1607 13730
rect 138 13648 172 13682
rect 231 13600 1607 13634
rect 1666 13552 1700 13586
rect 231 13504 1607 13538
rect 138 13456 172 13490
rect 231 13408 1607 13442
rect 1666 13360 1700 13394
rect 231 13312 1607 13346
rect 138 13264 172 13298
rect 231 13216 1607 13250
rect 1666 13168 1700 13202
rect 231 13120 1607 13154
rect 138 13072 172 13106
rect 231 13024 1607 13058
rect 1666 12976 1700 13010
rect 231 12928 1607 12962
rect 138 12880 172 12914
rect 231 12832 1607 12866
rect 1666 12784 1700 12818
rect 231 12736 1607 12770
rect 138 12688 172 12722
rect 231 12640 1607 12674
rect 1666 12592 1700 12626
rect 231 12544 1607 12578
rect 138 12496 172 12530
rect 231 12448 1607 12482
rect 1666 12400 1700 12434
rect 231 12352 1607 12386
rect 138 12304 172 12338
rect 231 12256 1607 12290
rect 1666 12208 1700 12242
rect 231 12160 1607 12194
rect 138 12112 172 12146
rect 231 12064 1607 12098
rect 1666 12016 1700 12050
rect 231 11968 1607 12002
rect 138 11920 172 11954
rect 231 11872 1607 11906
rect 1666 11824 1700 11858
rect 231 11776 1607 11810
rect 138 11728 172 11762
rect 231 11680 1607 11714
rect 1666 11632 1700 11666
rect 231 11584 1607 11618
rect 138 11536 172 11570
rect 231 11488 1607 11522
rect 1666 11440 1700 11474
rect 231 11392 1607 11426
rect 138 11344 172 11378
rect 231 11296 1607 11330
rect 1666 11248 1700 11282
rect 231 11200 1607 11234
rect 138 11152 172 11186
rect 231 11104 1607 11138
rect 1666 11056 1700 11090
rect 231 11008 1607 11042
rect 138 10960 172 10994
rect 231 10912 1607 10946
rect 1666 10864 1700 10898
rect 231 10816 1607 10850
rect 138 10768 172 10802
rect 231 10720 1607 10754
rect 1666 10672 1700 10706
rect 231 10624 1607 10658
rect 138 10576 172 10610
rect 231 10528 1607 10562
rect 1666 10480 1700 10514
rect 231 10432 1607 10466
rect 138 10384 172 10418
rect 231 10336 1607 10370
rect 1666 10288 1700 10322
rect 231 10240 1607 10274
rect 138 10192 172 10226
rect 231 10144 1607 10178
rect 1666 10096 1700 10130
rect 231 10048 1607 10082
rect 138 10000 172 10034
rect 231 9952 1607 9986
rect 1666 9904 1700 9938
rect 231 9856 1607 9890
rect 138 9808 172 9842
rect 231 9760 1607 9794
rect 1666 9712 1700 9746
rect 231 9664 1607 9698
rect 138 9616 172 9650
rect 231 9568 1607 9602
rect 1666 9520 1700 9554
rect 231 9472 1607 9506
rect 138 9424 172 9458
rect 231 9376 1607 9410
rect 1666 9328 1700 9362
rect 231 9280 1607 9314
rect 138 9232 172 9266
rect 231 9184 1607 9218
rect 1666 9136 1700 9170
rect 231 9088 1607 9122
rect 138 9040 172 9074
rect 231 8992 1607 9026
rect 1666 8944 1700 8978
rect 231 8896 1607 8930
rect 138 8848 172 8882
rect 231 8800 1607 8834
rect 1666 8752 1700 8786
rect 231 8704 1607 8738
rect 138 8656 172 8690
rect 231 8608 1607 8642
rect 1666 8560 1700 8594
rect 231 8512 1607 8546
rect 138 8464 172 8498
rect 231 8416 1607 8450
rect 1666 8368 1700 8402
rect 231 8320 1607 8354
rect 138 8272 172 8306
rect 231 8224 1607 8258
rect 1666 8176 1700 8210
rect 231 8128 1607 8162
rect 138 8080 172 8114
rect 231 8032 1607 8066
rect 1666 7984 1700 8018
rect 231 7936 1607 7970
rect 138 7888 172 7922
rect 231 7840 1607 7874
rect 1666 7792 1700 7826
rect 231 7744 1607 7778
rect 138 7696 172 7730
rect 231 7648 1607 7682
rect 1666 7600 1700 7634
rect 231 7552 1607 7586
rect 138 7504 172 7538
rect 231 7456 1607 7490
rect 1666 7408 1700 7442
rect 231 7360 1607 7394
rect 138 7312 172 7346
rect 231 7264 1607 7298
rect 1666 7216 1700 7250
rect 231 7168 1607 7202
rect 138 7120 172 7154
rect 231 7072 1607 7106
rect 1666 7024 1700 7058
rect 231 6976 1607 7010
rect 138 6928 172 6962
rect 231 6880 1607 6914
rect 1666 6832 1700 6866
rect 231 6784 1607 6818
rect 138 6736 172 6770
rect 231 6688 1607 6722
rect 1666 6640 1700 6674
rect 231 6592 1607 6626
rect 138 6544 172 6578
rect 231 6496 1607 6530
rect 1666 6448 1700 6482
rect 231 6400 1607 6434
rect 138 6352 172 6386
rect 231 6304 1607 6338
rect 1666 6256 1700 6290
rect 231 6208 1607 6242
rect 138 6160 172 6194
rect 231 6112 1607 6146
rect 1666 6064 1700 6098
rect 231 6016 1607 6050
rect 138 5968 172 6002
rect 231 5920 1607 5954
rect 1666 5872 1700 5906
rect 231 5824 1607 5858
rect 138 5776 172 5810
rect 231 5728 1607 5762
rect 1666 5680 1700 5714
rect 231 5632 1607 5666
rect 138 5584 172 5618
rect 231 5536 1607 5570
rect 1666 5488 1700 5522
rect 231 5440 1607 5474
rect 138 5392 172 5426
rect 231 5344 1607 5378
rect 1666 5296 1700 5330
rect 231 5248 1607 5282
rect 138 5200 172 5234
rect 231 5152 1607 5186
rect 1666 5104 1700 5138
rect 231 5056 1607 5090
rect 138 5008 172 5042
rect 231 4960 1607 4994
rect 1666 4912 1700 4946
rect 231 4864 1607 4898
rect 138 4816 172 4850
rect 231 4768 1607 4802
rect 1666 4720 1700 4754
rect 231 4672 1607 4706
rect 138 4624 172 4658
rect 231 4576 1607 4610
rect 1666 4528 1700 4562
rect 231 4480 1607 4514
rect 138 4432 172 4466
rect 231 4384 1607 4418
rect 1666 4336 1700 4370
rect 231 4288 1607 4322
rect 138 4240 172 4274
rect 231 4192 1607 4226
rect 1666 4144 1700 4178
rect 231 4096 1607 4130
rect 138 4048 172 4082
rect 231 4000 1607 4034
rect 1666 3952 1700 3986
rect 231 3904 1607 3938
rect 138 3856 172 3890
rect 231 3808 1607 3842
rect 1666 3760 1700 3794
rect 231 3712 1607 3746
rect 138 3664 172 3698
rect 231 3616 1607 3650
rect 1666 3568 1700 3602
rect 231 3520 1607 3554
rect 138 3472 172 3506
rect 231 3424 1607 3458
rect 1666 3376 1700 3410
rect 231 3328 1607 3362
rect 138 3280 172 3314
rect 231 3232 1607 3266
rect 1666 3184 1700 3218
rect 231 3136 1607 3170
rect 138 3088 172 3122
rect 231 3040 1607 3074
rect 1666 2992 1700 3026
rect 231 2944 1607 2978
rect 138 2896 172 2930
rect 231 2848 1607 2882
rect 1666 2800 1700 2834
rect 231 2752 1607 2786
rect 138 2704 172 2738
rect 231 2656 1607 2690
rect 1666 2608 1700 2642
rect 231 2560 1607 2594
rect 138 2512 172 2546
rect 231 2464 1607 2498
rect 1666 2416 1700 2450
rect 231 2368 1607 2402
rect 138 2320 172 2354
rect 231 2272 1607 2306
rect 1666 2224 1700 2258
rect 231 2176 1607 2210
rect 138 2128 172 2162
rect 231 2080 1607 2114
rect 1666 2032 1700 2066
rect 231 1984 1607 2018
rect 138 1936 172 1970
rect 231 1888 1607 1922
rect 1666 1840 1700 1874
rect 231 1792 1607 1826
rect 138 1744 172 1778
rect 231 1696 1607 1730
rect 1666 1648 1700 1682
rect 231 1600 1607 1634
rect 138 1552 172 1586
rect 231 1504 1607 1538
rect 1666 1456 1700 1490
rect 231 1408 1607 1442
rect 138 1360 172 1394
rect 231 1312 1607 1346
rect 1666 1264 1700 1298
rect 231 1216 1607 1250
rect 138 1168 172 1202
rect 231 1120 1607 1154
rect 1666 1072 1700 1106
rect 231 1024 1607 1058
rect 138 976 172 1010
rect 231 928 1607 962
rect 1666 880 1700 914
rect 231 832 1607 866
rect 138 784 172 818
rect 231 736 1607 770
rect 1666 688 1700 722
rect 231 640 1607 674
<< metal1 >>
rect 122 22286 1716 22304
rect 122 22222 132 22286
rect 1706 22222 1716 22286
rect 122 22204 1716 22222
rect 132 21746 178 22204
rect 316 21934 894 21938
rect 316 21932 352 21934
rect 858 21932 894 21934
rect 316 21868 328 21932
rect 882 21868 894 21932
rect 316 21862 894 21868
rect 342 21800 352 21810
rect 219 21794 352 21800
rect 858 21800 868 21810
rect 858 21794 1619 21800
rect 219 21760 231 21794
rect 1607 21760 1619 21794
rect 219 21754 352 21760
rect 132 21712 138 21746
rect 172 21712 178 21746
rect 342 21744 352 21754
rect 858 21754 1619 21760
rect 858 21744 868 21754
rect 132 21554 178 21712
rect 970 21704 980 21714
rect 219 21698 980 21704
rect 1490 21704 1500 21714
rect 1490 21698 1619 21704
rect 219 21664 231 21698
rect 1607 21664 1619 21698
rect 219 21658 980 21664
rect 970 21648 980 21658
rect 1490 21658 1619 21664
rect 1490 21648 1500 21658
rect 1660 21650 1706 22204
rect 342 21608 352 21618
rect 219 21602 352 21608
rect 858 21608 868 21618
rect 1660 21616 1666 21650
rect 1700 21616 1706 21650
rect 858 21602 1619 21608
rect 219 21568 231 21602
rect 1607 21568 1619 21602
rect 219 21562 352 21568
rect 132 21520 138 21554
rect 172 21520 178 21554
rect 342 21552 352 21562
rect 858 21562 1619 21568
rect 858 21552 868 21562
rect 132 21362 178 21520
rect 970 21512 980 21522
rect 219 21506 980 21512
rect 1490 21512 1500 21522
rect 1490 21506 1619 21512
rect 219 21472 231 21506
rect 1607 21472 1619 21506
rect 219 21466 980 21472
rect 970 21456 980 21466
rect 1490 21466 1619 21472
rect 1490 21456 1500 21466
rect 1660 21458 1706 21616
rect 342 21416 352 21426
rect 219 21410 352 21416
rect 858 21416 868 21426
rect 1660 21424 1666 21458
rect 1700 21424 1706 21458
rect 858 21410 1619 21416
rect 219 21376 231 21410
rect 1607 21376 1619 21410
rect 219 21370 352 21376
rect 132 21328 138 21362
rect 172 21328 178 21362
rect 342 21360 352 21370
rect 858 21370 1619 21376
rect 858 21360 868 21370
rect 132 21170 178 21328
rect 970 21320 980 21330
rect 219 21314 980 21320
rect 1490 21320 1500 21330
rect 1490 21314 1619 21320
rect 219 21280 231 21314
rect 1607 21280 1619 21314
rect 219 21274 980 21280
rect 970 21264 980 21274
rect 1490 21274 1619 21280
rect 1490 21264 1500 21274
rect 1660 21266 1706 21424
rect 342 21224 352 21234
rect 219 21218 352 21224
rect 858 21224 868 21234
rect 1660 21232 1666 21266
rect 1700 21232 1706 21266
rect 858 21218 1619 21224
rect 219 21184 231 21218
rect 1607 21184 1619 21218
rect 219 21178 352 21184
rect 132 21136 138 21170
rect 172 21136 178 21170
rect 342 21168 352 21178
rect 858 21178 1619 21184
rect 858 21168 868 21178
rect 132 20978 178 21136
rect 970 21128 980 21138
rect 219 21122 980 21128
rect 1490 21128 1500 21138
rect 1490 21122 1619 21128
rect 219 21088 231 21122
rect 1607 21088 1619 21122
rect 219 21082 980 21088
rect 970 21072 980 21082
rect 1490 21082 1619 21088
rect 1490 21072 1500 21082
rect 1660 21074 1706 21232
rect 342 21032 352 21042
rect 219 21026 352 21032
rect 858 21032 868 21042
rect 1660 21040 1666 21074
rect 1700 21040 1706 21074
rect 858 21026 1619 21032
rect 219 20992 231 21026
rect 1607 20992 1619 21026
rect 219 20986 352 20992
rect 132 20944 138 20978
rect 172 20944 178 20978
rect 342 20976 352 20986
rect 858 20986 1619 20992
rect 858 20976 868 20986
rect 132 20786 178 20944
rect 970 20936 980 20946
rect 219 20930 980 20936
rect 1490 20936 1500 20946
rect 1490 20930 1619 20936
rect 219 20896 231 20930
rect 1607 20896 1619 20930
rect 219 20890 980 20896
rect 970 20880 980 20890
rect 1490 20890 1619 20896
rect 1490 20880 1500 20890
rect 1660 20882 1706 21040
rect 342 20840 352 20850
rect 219 20834 352 20840
rect 858 20840 868 20850
rect 1660 20848 1666 20882
rect 1700 20848 1706 20882
rect 858 20834 1619 20840
rect 219 20800 231 20834
rect 1607 20800 1619 20834
rect 219 20794 352 20800
rect 132 20752 138 20786
rect 172 20752 178 20786
rect 342 20784 352 20794
rect 858 20794 1619 20800
rect 858 20784 868 20794
rect 132 20594 178 20752
rect 970 20744 980 20754
rect 219 20738 980 20744
rect 1490 20744 1500 20754
rect 1490 20738 1619 20744
rect 219 20704 231 20738
rect 1607 20704 1619 20738
rect 219 20698 980 20704
rect 970 20688 980 20698
rect 1490 20698 1619 20704
rect 1490 20688 1500 20698
rect 1660 20690 1706 20848
rect 342 20648 352 20658
rect 219 20642 352 20648
rect 858 20648 868 20658
rect 1660 20656 1666 20690
rect 1700 20656 1706 20690
rect 858 20642 1619 20648
rect 219 20608 231 20642
rect 1607 20608 1619 20642
rect 219 20602 352 20608
rect 132 20560 138 20594
rect 172 20560 178 20594
rect 342 20592 352 20602
rect 858 20602 1619 20608
rect 858 20592 868 20602
rect 132 20402 178 20560
rect 970 20552 980 20562
rect 219 20546 980 20552
rect 1490 20552 1500 20562
rect 1490 20546 1619 20552
rect 219 20512 231 20546
rect 1607 20512 1619 20546
rect 219 20506 980 20512
rect 970 20496 980 20506
rect 1490 20506 1619 20512
rect 1490 20496 1500 20506
rect 1660 20498 1706 20656
rect 342 20456 352 20466
rect 219 20450 352 20456
rect 858 20456 868 20466
rect 1660 20464 1666 20498
rect 1700 20464 1706 20498
rect 858 20450 1619 20456
rect 219 20416 231 20450
rect 1607 20416 1619 20450
rect 219 20410 352 20416
rect 132 20368 138 20402
rect 172 20368 178 20402
rect 342 20400 352 20410
rect 858 20410 1619 20416
rect 858 20400 868 20410
rect 132 20210 178 20368
rect 970 20360 980 20370
rect 219 20354 980 20360
rect 1490 20360 1500 20370
rect 1490 20354 1619 20360
rect 219 20320 231 20354
rect 1607 20320 1619 20354
rect 219 20314 980 20320
rect 970 20304 980 20314
rect 1490 20314 1619 20320
rect 1490 20304 1500 20314
rect 1660 20306 1706 20464
rect 342 20264 352 20274
rect 219 20258 352 20264
rect 858 20264 868 20274
rect 1660 20272 1666 20306
rect 1700 20272 1706 20306
rect 858 20258 1619 20264
rect 219 20224 231 20258
rect 1607 20224 1619 20258
rect 219 20218 352 20224
rect 132 20176 138 20210
rect 172 20176 178 20210
rect 342 20208 352 20218
rect 858 20218 1619 20224
rect 858 20208 868 20218
rect 132 20018 178 20176
rect 970 20168 980 20178
rect 219 20162 980 20168
rect 1490 20168 1500 20178
rect 1490 20162 1619 20168
rect 219 20128 231 20162
rect 1607 20128 1619 20162
rect 219 20122 980 20128
rect 970 20112 980 20122
rect 1490 20122 1619 20128
rect 1490 20112 1500 20122
rect 1660 20114 1706 20272
rect 342 20072 352 20082
rect 219 20066 352 20072
rect 858 20072 868 20082
rect 1660 20080 1666 20114
rect 1700 20080 1706 20114
rect 858 20066 1619 20072
rect 219 20032 231 20066
rect 1607 20032 1619 20066
rect 219 20026 352 20032
rect 132 19984 138 20018
rect 172 19984 178 20018
rect 342 20016 352 20026
rect 858 20026 1619 20032
rect 858 20016 868 20026
rect 132 19826 178 19984
rect 970 19976 980 19986
rect 219 19970 980 19976
rect 1490 19976 1500 19986
rect 1490 19970 1619 19976
rect 219 19936 231 19970
rect 1607 19936 1619 19970
rect 219 19930 980 19936
rect 970 19920 980 19930
rect 1490 19930 1619 19936
rect 1490 19920 1500 19930
rect 1660 19922 1706 20080
rect 342 19880 352 19890
rect 219 19874 352 19880
rect 858 19880 868 19890
rect 1660 19888 1666 19922
rect 1700 19888 1706 19922
rect 858 19874 1619 19880
rect 219 19840 231 19874
rect 1607 19840 1619 19874
rect 219 19834 352 19840
rect 132 19792 138 19826
rect 172 19792 178 19826
rect 342 19824 352 19834
rect 858 19834 1619 19840
rect 858 19824 868 19834
rect 132 19634 178 19792
rect 970 19784 980 19794
rect 219 19778 980 19784
rect 1490 19784 1500 19794
rect 1490 19778 1619 19784
rect 219 19744 231 19778
rect 1607 19744 1619 19778
rect 219 19738 980 19744
rect 970 19728 980 19738
rect 1490 19738 1619 19744
rect 1490 19728 1500 19738
rect 1660 19730 1706 19888
rect 342 19688 352 19698
rect 219 19682 352 19688
rect 858 19688 868 19698
rect 1660 19696 1666 19730
rect 1700 19696 1706 19730
rect 858 19682 1619 19688
rect 219 19648 231 19682
rect 1607 19648 1619 19682
rect 219 19642 352 19648
rect 132 19600 138 19634
rect 172 19600 178 19634
rect 342 19632 352 19642
rect 858 19642 1619 19648
rect 858 19632 868 19642
rect 132 19442 178 19600
rect 970 19592 980 19602
rect 219 19586 980 19592
rect 1490 19592 1500 19602
rect 1490 19586 1619 19592
rect 219 19552 231 19586
rect 1607 19552 1619 19586
rect 219 19546 980 19552
rect 970 19536 980 19546
rect 1490 19546 1619 19552
rect 1490 19536 1500 19546
rect 1660 19538 1706 19696
rect 342 19496 352 19506
rect 219 19490 352 19496
rect 858 19496 868 19506
rect 1660 19504 1666 19538
rect 1700 19504 1706 19538
rect 858 19490 1619 19496
rect 219 19456 231 19490
rect 1607 19456 1619 19490
rect 219 19450 352 19456
rect 132 19408 138 19442
rect 172 19408 178 19442
rect 342 19440 352 19450
rect 858 19450 1619 19456
rect 858 19440 868 19450
rect 132 19250 178 19408
rect 970 19400 980 19410
rect 219 19394 980 19400
rect 1490 19400 1500 19410
rect 1490 19394 1619 19400
rect 219 19360 231 19394
rect 1607 19360 1619 19394
rect 219 19354 980 19360
rect 970 19344 980 19354
rect 1490 19354 1619 19360
rect 1490 19344 1500 19354
rect 1660 19346 1706 19504
rect 342 19304 352 19314
rect 219 19298 352 19304
rect 858 19304 868 19314
rect 1660 19312 1666 19346
rect 1700 19312 1706 19346
rect 858 19298 1619 19304
rect 219 19264 231 19298
rect 1607 19264 1619 19298
rect 219 19258 352 19264
rect 132 19216 138 19250
rect 172 19216 178 19250
rect 342 19248 352 19258
rect 858 19258 1619 19264
rect 858 19248 868 19258
rect 132 19058 178 19216
rect 970 19208 980 19218
rect 219 19202 980 19208
rect 1490 19208 1500 19218
rect 1490 19202 1619 19208
rect 219 19168 231 19202
rect 1607 19168 1619 19202
rect 219 19162 980 19168
rect 970 19152 980 19162
rect 1490 19162 1619 19168
rect 1490 19152 1500 19162
rect 1660 19154 1706 19312
rect 342 19112 352 19122
rect 219 19106 352 19112
rect 858 19112 868 19122
rect 1660 19120 1666 19154
rect 1700 19120 1706 19154
rect 858 19106 1619 19112
rect 219 19072 231 19106
rect 1607 19072 1619 19106
rect 219 19066 352 19072
rect 132 19024 138 19058
rect 172 19024 178 19058
rect 342 19056 352 19066
rect 858 19066 1619 19072
rect 858 19056 868 19066
rect 132 18866 178 19024
rect 970 19016 980 19026
rect 219 19010 980 19016
rect 1490 19016 1500 19026
rect 1490 19010 1619 19016
rect 219 18976 231 19010
rect 1607 18976 1619 19010
rect 219 18970 980 18976
rect 970 18960 980 18970
rect 1490 18970 1619 18976
rect 1490 18960 1500 18970
rect 1660 18962 1706 19120
rect 342 18920 352 18930
rect 219 18914 352 18920
rect 858 18920 868 18930
rect 1660 18928 1666 18962
rect 1700 18928 1706 18962
rect 858 18914 1619 18920
rect 219 18880 231 18914
rect 1607 18880 1619 18914
rect 219 18874 352 18880
rect 132 18832 138 18866
rect 172 18832 178 18866
rect 342 18864 352 18874
rect 858 18874 1619 18880
rect 858 18864 868 18874
rect 132 18674 178 18832
rect 970 18824 980 18834
rect 219 18818 980 18824
rect 1490 18824 1500 18834
rect 1490 18818 1619 18824
rect 219 18784 231 18818
rect 1607 18784 1619 18818
rect 219 18778 980 18784
rect 970 18768 980 18778
rect 1490 18778 1619 18784
rect 1490 18768 1500 18778
rect 1660 18770 1706 18928
rect 342 18728 352 18738
rect 219 18722 352 18728
rect 858 18728 868 18738
rect 1660 18736 1666 18770
rect 1700 18736 1706 18770
rect 858 18722 1619 18728
rect 219 18688 231 18722
rect 1607 18688 1619 18722
rect 219 18682 352 18688
rect 132 18640 138 18674
rect 172 18640 178 18674
rect 342 18672 352 18682
rect 858 18682 1619 18688
rect 858 18672 868 18682
rect 132 18482 178 18640
rect 970 18632 980 18642
rect 219 18626 980 18632
rect 1490 18632 1500 18642
rect 1490 18626 1619 18632
rect 219 18592 231 18626
rect 1607 18592 1619 18626
rect 219 18586 980 18592
rect 970 18576 980 18586
rect 1490 18586 1619 18592
rect 1490 18576 1500 18586
rect 1660 18578 1706 18736
rect 342 18536 352 18546
rect 219 18530 352 18536
rect 858 18536 868 18546
rect 1660 18544 1666 18578
rect 1700 18544 1706 18578
rect 858 18530 1619 18536
rect 219 18496 231 18530
rect 1607 18496 1619 18530
rect 219 18490 352 18496
rect 132 18448 138 18482
rect 172 18448 178 18482
rect 342 18480 352 18490
rect 858 18490 1619 18496
rect 858 18480 868 18490
rect 132 18290 178 18448
rect 970 18440 980 18450
rect 219 18434 980 18440
rect 1490 18440 1500 18450
rect 1490 18434 1619 18440
rect 219 18400 231 18434
rect 1607 18400 1619 18434
rect 219 18394 980 18400
rect 970 18384 980 18394
rect 1490 18394 1619 18400
rect 1490 18384 1500 18394
rect 1660 18386 1706 18544
rect 342 18344 352 18354
rect 219 18338 352 18344
rect 858 18344 868 18354
rect 1660 18352 1666 18386
rect 1700 18352 1706 18386
rect 858 18338 1619 18344
rect 219 18304 231 18338
rect 1607 18304 1619 18338
rect 219 18298 352 18304
rect 132 18256 138 18290
rect 172 18256 178 18290
rect 342 18288 352 18298
rect 858 18298 1619 18304
rect 858 18288 868 18298
rect 132 18098 178 18256
rect 970 18248 980 18258
rect 219 18242 980 18248
rect 1490 18248 1500 18258
rect 1490 18242 1619 18248
rect 219 18208 231 18242
rect 1607 18208 1619 18242
rect 219 18202 980 18208
rect 970 18192 980 18202
rect 1490 18202 1619 18208
rect 1490 18192 1500 18202
rect 1660 18194 1706 18352
rect 342 18152 352 18162
rect 219 18146 352 18152
rect 858 18152 868 18162
rect 1660 18160 1666 18194
rect 1700 18160 1706 18194
rect 858 18146 1619 18152
rect 219 18112 231 18146
rect 1607 18112 1619 18146
rect 219 18106 352 18112
rect 132 18064 138 18098
rect 172 18064 178 18098
rect 342 18096 352 18106
rect 858 18106 1619 18112
rect 858 18096 868 18106
rect 132 17906 178 18064
rect 970 18056 980 18066
rect 219 18050 980 18056
rect 1490 18056 1500 18066
rect 1490 18050 1619 18056
rect 219 18016 231 18050
rect 1607 18016 1619 18050
rect 219 18010 980 18016
rect 970 18000 980 18010
rect 1490 18010 1619 18016
rect 1490 18000 1500 18010
rect 1660 18002 1706 18160
rect 342 17960 352 17970
rect 219 17954 352 17960
rect 858 17960 868 17970
rect 1660 17968 1666 18002
rect 1700 17968 1706 18002
rect 858 17954 1619 17960
rect 219 17920 231 17954
rect 1607 17920 1619 17954
rect 219 17914 352 17920
rect 132 17872 138 17906
rect 172 17872 178 17906
rect 342 17904 352 17914
rect 858 17914 1619 17920
rect 858 17904 868 17914
rect 132 17714 178 17872
rect 970 17864 980 17874
rect 219 17858 980 17864
rect 1490 17864 1500 17874
rect 1490 17858 1619 17864
rect 219 17824 231 17858
rect 1607 17824 1619 17858
rect 219 17818 980 17824
rect 970 17808 980 17818
rect 1490 17818 1619 17824
rect 1490 17808 1500 17818
rect 1660 17810 1706 17968
rect 342 17768 352 17778
rect 219 17762 352 17768
rect 858 17768 868 17778
rect 1660 17776 1666 17810
rect 1700 17776 1706 17810
rect 858 17762 1619 17768
rect 219 17728 231 17762
rect 1607 17728 1619 17762
rect 219 17722 352 17728
rect 132 17680 138 17714
rect 172 17680 178 17714
rect 342 17712 352 17722
rect 858 17722 1619 17728
rect 858 17712 868 17722
rect 132 17522 178 17680
rect 970 17672 980 17682
rect 219 17666 980 17672
rect 1490 17672 1500 17682
rect 1490 17666 1619 17672
rect 219 17632 231 17666
rect 1607 17632 1619 17666
rect 219 17626 980 17632
rect 970 17616 980 17626
rect 1490 17626 1619 17632
rect 1490 17616 1500 17626
rect 1660 17618 1706 17776
rect 342 17576 352 17586
rect 219 17570 352 17576
rect 858 17576 868 17586
rect 1660 17584 1666 17618
rect 1700 17584 1706 17618
rect 858 17570 1619 17576
rect 219 17536 231 17570
rect 1607 17536 1619 17570
rect 219 17530 352 17536
rect 132 17488 138 17522
rect 172 17488 178 17522
rect 342 17520 352 17530
rect 858 17530 1619 17536
rect 858 17520 868 17530
rect 132 17330 178 17488
rect 970 17480 980 17490
rect 219 17474 980 17480
rect 1490 17480 1500 17490
rect 1490 17474 1619 17480
rect 219 17440 231 17474
rect 1607 17440 1619 17474
rect 219 17434 980 17440
rect 970 17424 980 17434
rect 1490 17434 1619 17440
rect 1490 17424 1500 17434
rect 1660 17426 1706 17584
rect 342 17384 352 17394
rect 219 17378 352 17384
rect 858 17384 868 17394
rect 1660 17392 1666 17426
rect 1700 17392 1706 17426
rect 858 17378 1619 17384
rect 219 17344 231 17378
rect 1607 17344 1619 17378
rect 219 17338 352 17344
rect 132 17296 138 17330
rect 172 17296 178 17330
rect 342 17328 352 17338
rect 858 17338 1619 17344
rect 858 17328 868 17338
rect 132 17138 178 17296
rect 970 17288 980 17298
rect 219 17282 980 17288
rect 1490 17288 1500 17298
rect 1490 17282 1619 17288
rect 219 17248 231 17282
rect 1607 17248 1619 17282
rect 219 17242 980 17248
rect 970 17232 980 17242
rect 1490 17242 1619 17248
rect 1490 17232 1500 17242
rect 1660 17234 1706 17392
rect 342 17192 352 17202
rect 219 17186 352 17192
rect 858 17192 868 17202
rect 1660 17200 1666 17234
rect 1700 17200 1706 17234
rect 858 17186 1619 17192
rect 219 17152 231 17186
rect 1607 17152 1619 17186
rect 219 17146 352 17152
rect 132 17104 138 17138
rect 172 17104 178 17138
rect 342 17136 352 17146
rect 858 17146 1619 17152
rect 858 17136 868 17146
rect 132 16946 178 17104
rect 970 17096 980 17106
rect 219 17090 980 17096
rect 1490 17096 1500 17106
rect 1490 17090 1619 17096
rect 219 17056 231 17090
rect 1607 17056 1619 17090
rect 219 17050 980 17056
rect 970 17040 980 17050
rect 1490 17050 1619 17056
rect 1490 17040 1500 17050
rect 1660 17042 1706 17200
rect 342 17000 352 17010
rect 219 16994 352 17000
rect 858 17000 868 17010
rect 1660 17008 1666 17042
rect 1700 17008 1706 17042
rect 858 16994 1619 17000
rect 219 16960 231 16994
rect 1607 16960 1619 16994
rect 219 16954 352 16960
rect 132 16912 138 16946
rect 172 16912 178 16946
rect 342 16944 352 16954
rect 858 16954 1619 16960
rect 858 16944 868 16954
rect 132 16754 178 16912
rect 970 16904 980 16914
rect 219 16898 980 16904
rect 1490 16904 1500 16914
rect 1490 16898 1619 16904
rect 219 16864 231 16898
rect 1607 16864 1619 16898
rect 219 16858 980 16864
rect 970 16848 980 16858
rect 1490 16858 1619 16864
rect 1490 16848 1500 16858
rect 1660 16850 1706 17008
rect 342 16808 352 16818
rect 219 16802 352 16808
rect 858 16808 868 16818
rect 1660 16816 1666 16850
rect 1700 16816 1706 16850
rect 858 16802 1619 16808
rect 219 16768 231 16802
rect 1607 16768 1619 16802
rect 219 16762 352 16768
rect 132 16720 138 16754
rect 172 16720 178 16754
rect 342 16752 352 16762
rect 858 16762 1619 16768
rect 858 16752 868 16762
rect 132 16562 178 16720
rect 970 16712 980 16722
rect 219 16706 980 16712
rect 1490 16712 1500 16722
rect 1490 16706 1619 16712
rect 219 16672 231 16706
rect 1607 16672 1619 16706
rect 219 16666 980 16672
rect 970 16656 980 16666
rect 1490 16666 1619 16672
rect 1490 16656 1500 16666
rect 1660 16658 1706 16816
rect 342 16616 352 16626
rect 219 16610 352 16616
rect 858 16616 868 16626
rect 1660 16624 1666 16658
rect 1700 16624 1706 16658
rect 858 16610 1619 16616
rect 219 16576 231 16610
rect 1607 16576 1619 16610
rect 219 16570 352 16576
rect 132 16528 138 16562
rect 172 16528 178 16562
rect 342 16560 352 16570
rect 858 16570 1619 16576
rect 858 16560 868 16570
rect 132 16370 178 16528
rect 970 16520 980 16530
rect 219 16514 980 16520
rect 1490 16520 1500 16530
rect 1490 16514 1619 16520
rect 219 16480 231 16514
rect 1607 16480 1619 16514
rect 219 16474 980 16480
rect 970 16464 980 16474
rect 1490 16474 1619 16480
rect 1490 16464 1500 16474
rect 1660 16466 1706 16624
rect 342 16424 352 16434
rect 219 16418 352 16424
rect 858 16424 868 16434
rect 1660 16432 1666 16466
rect 1700 16432 1706 16466
rect 858 16418 1619 16424
rect 219 16384 231 16418
rect 1607 16384 1619 16418
rect 219 16378 352 16384
rect 132 16336 138 16370
rect 172 16336 178 16370
rect 342 16368 352 16378
rect 858 16378 1619 16384
rect 858 16368 868 16378
rect 132 16178 178 16336
rect 970 16328 980 16338
rect 219 16322 980 16328
rect 1490 16328 1500 16338
rect 1490 16322 1619 16328
rect 219 16288 231 16322
rect 1607 16288 1619 16322
rect 219 16282 980 16288
rect 970 16272 980 16282
rect 1490 16282 1619 16288
rect 1490 16272 1500 16282
rect 1660 16274 1706 16432
rect 342 16232 352 16242
rect 219 16226 352 16232
rect 858 16232 868 16242
rect 1660 16240 1666 16274
rect 1700 16240 1706 16274
rect 858 16226 1619 16232
rect 219 16192 231 16226
rect 1607 16192 1619 16226
rect 219 16186 352 16192
rect 132 16144 138 16178
rect 172 16144 178 16178
rect 342 16176 352 16186
rect 858 16186 1619 16192
rect 858 16176 868 16186
rect 132 15986 178 16144
rect 970 16136 980 16146
rect 219 16130 980 16136
rect 1490 16136 1500 16146
rect 1490 16130 1619 16136
rect 219 16096 231 16130
rect 1607 16096 1619 16130
rect 219 16090 980 16096
rect 970 16080 980 16090
rect 1490 16090 1619 16096
rect 1490 16080 1500 16090
rect 1660 16082 1706 16240
rect 342 16040 352 16050
rect 219 16034 352 16040
rect 858 16040 868 16050
rect 1660 16048 1666 16082
rect 1700 16048 1706 16082
rect 858 16034 1619 16040
rect 219 16000 231 16034
rect 1607 16000 1619 16034
rect 219 15994 352 16000
rect 132 15952 138 15986
rect 172 15952 178 15986
rect 342 15984 352 15994
rect 858 15994 1619 16000
rect 858 15984 868 15994
rect 132 15794 178 15952
rect 970 15944 980 15954
rect 219 15938 980 15944
rect 1490 15944 1500 15954
rect 1490 15938 1619 15944
rect 219 15904 231 15938
rect 1607 15904 1619 15938
rect 219 15898 980 15904
rect 970 15888 980 15898
rect 1490 15898 1619 15904
rect 1490 15888 1500 15898
rect 1660 15890 1706 16048
rect 342 15848 352 15858
rect 219 15842 352 15848
rect 858 15848 868 15858
rect 1660 15856 1666 15890
rect 1700 15856 1706 15890
rect 858 15842 1619 15848
rect 219 15808 231 15842
rect 1607 15808 1619 15842
rect 219 15802 352 15808
rect 132 15760 138 15794
rect 172 15760 178 15794
rect 342 15792 352 15802
rect 858 15802 1619 15808
rect 858 15792 868 15802
rect 132 15602 178 15760
rect 970 15752 980 15762
rect 219 15746 980 15752
rect 1490 15752 1500 15762
rect 1490 15746 1619 15752
rect 219 15712 231 15746
rect 1607 15712 1619 15746
rect 219 15706 980 15712
rect 970 15696 980 15706
rect 1490 15706 1619 15712
rect 1490 15696 1500 15706
rect 1660 15698 1706 15856
rect 342 15656 352 15666
rect 219 15650 352 15656
rect 858 15656 868 15666
rect 1660 15664 1666 15698
rect 1700 15664 1706 15698
rect 858 15650 1619 15656
rect 219 15616 231 15650
rect 1607 15616 1619 15650
rect 219 15610 352 15616
rect 132 15568 138 15602
rect 172 15568 178 15602
rect 342 15600 352 15610
rect 858 15610 1619 15616
rect 858 15600 868 15610
rect 132 15410 178 15568
rect 970 15560 980 15570
rect 219 15554 980 15560
rect 1490 15560 1500 15570
rect 1490 15554 1619 15560
rect 219 15520 231 15554
rect 1607 15520 1619 15554
rect 219 15514 980 15520
rect 970 15504 980 15514
rect 1490 15514 1619 15520
rect 1490 15504 1500 15514
rect 1660 15506 1706 15664
rect 342 15464 352 15474
rect 219 15458 352 15464
rect 858 15464 868 15474
rect 1660 15472 1666 15506
rect 1700 15472 1706 15506
rect 858 15458 1619 15464
rect 219 15424 231 15458
rect 1607 15424 1619 15458
rect 219 15418 352 15424
rect 132 15376 138 15410
rect 172 15376 178 15410
rect 342 15408 352 15418
rect 858 15418 1619 15424
rect 858 15408 868 15418
rect 132 15218 178 15376
rect 970 15368 980 15378
rect 219 15362 980 15368
rect 1490 15368 1500 15378
rect 1490 15362 1619 15368
rect 219 15328 231 15362
rect 1607 15328 1619 15362
rect 219 15322 980 15328
rect 970 15312 980 15322
rect 1490 15322 1619 15328
rect 1490 15312 1500 15322
rect 1660 15314 1706 15472
rect 342 15272 352 15282
rect 219 15266 352 15272
rect 858 15272 868 15282
rect 1660 15280 1666 15314
rect 1700 15280 1706 15314
rect 858 15266 1619 15272
rect 219 15232 231 15266
rect 1607 15232 1619 15266
rect 219 15226 352 15232
rect 132 15184 138 15218
rect 172 15184 178 15218
rect 342 15216 352 15226
rect 858 15226 1619 15232
rect 858 15216 868 15226
rect 132 15026 178 15184
rect 970 15176 980 15186
rect 219 15170 980 15176
rect 1490 15176 1500 15186
rect 1490 15170 1619 15176
rect 219 15136 231 15170
rect 1607 15136 1619 15170
rect 219 15130 980 15136
rect 970 15120 980 15130
rect 1490 15130 1619 15136
rect 1490 15120 1500 15130
rect 1660 15122 1706 15280
rect 342 15080 352 15090
rect 219 15074 352 15080
rect 858 15080 868 15090
rect 1660 15088 1666 15122
rect 1700 15088 1706 15122
rect 858 15074 1619 15080
rect 219 15040 231 15074
rect 1607 15040 1619 15074
rect 219 15034 352 15040
rect 132 14992 138 15026
rect 172 14992 178 15026
rect 342 15024 352 15034
rect 858 15034 1619 15040
rect 858 15024 868 15034
rect 132 14834 178 14992
rect 970 14984 980 14994
rect 219 14978 980 14984
rect 1490 14984 1500 14994
rect 1490 14978 1619 14984
rect 219 14944 231 14978
rect 1607 14944 1619 14978
rect 219 14938 980 14944
rect 970 14928 980 14938
rect 1490 14938 1619 14944
rect 1490 14928 1500 14938
rect 1660 14930 1706 15088
rect 342 14888 352 14898
rect 219 14882 352 14888
rect 858 14888 868 14898
rect 1660 14896 1666 14930
rect 1700 14896 1706 14930
rect 858 14882 1619 14888
rect 219 14848 231 14882
rect 1607 14848 1619 14882
rect 219 14842 352 14848
rect 132 14800 138 14834
rect 172 14800 178 14834
rect 342 14832 352 14842
rect 858 14842 1619 14848
rect 858 14832 868 14842
rect 132 14642 178 14800
rect 970 14792 980 14802
rect 219 14786 980 14792
rect 1490 14792 1500 14802
rect 1490 14786 1619 14792
rect 219 14752 231 14786
rect 1607 14752 1619 14786
rect 219 14746 980 14752
rect 970 14736 980 14746
rect 1490 14746 1619 14752
rect 1490 14736 1500 14746
rect 1660 14738 1706 14896
rect 342 14696 352 14706
rect 219 14690 352 14696
rect 858 14696 868 14706
rect 1660 14704 1666 14738
rect 1700 14704 1706 14738
rect 858 14690 1619 14696
rect 219 14656 231 14690
rect 1607 14656 1619 14690
rect 219 14650 352 14656
rect 132 14608 138 14642
rect 172 14608 178 14642
rect 342 14640 352 14650
rect 858 14650 1619 14656
rect 858 14640 868 14650
rect 132 14450 178 14608
rect 970 14600 980 14610
rect 219 14594 980 14600
rect 1490 14600 1500 14610
rect 1490 14594 1619 14600
rect 219 14560 231 14594
rect 1607 14560 1619 14594
rect 219 14554 980 14560
rect 970 14544 980 14554
rect 1490 14554 1619 14560
rect 1490 14544 1500 14554
rect 1660 14546 1706 14704
rect 342 14504 352 14514
rect 219 14498 352 14504
rect 858 14504 868 14514
rect 1660 14512 1666 14546
rect 1700 14512 1706 14546
rect 858 14498 1619 14504
rect 219 14464 231 14498
rect 1607 14464 1619 14498
rect 219 14458 352 14464
rect 132 14416 138 14450
rect 172 14416 178 14450
rect 342 14448 352 14458
rect 858 14458 1619 14464
rect 858 14448 868 14458
rect 132 14258 178 14416
rect 970 14408 980 14418
rect 219 14402 980 14408
rect 1490 14408 1500 14418
rect 1490 14402 1619 14408
rect 219 14368 231 14402
rect 1607 14368 1619 14402
rect 219 14362 980 14368
rect 970 14352 980 14362
rect 1490 14362 1619 14368
rect 1490 14352 1500 14362
rect 1660 14354 1706 14512
rect 342 14312 352 14322
rect 219 14306 352 14312
rect 858 14312 868 14322
rect 1660 14320 1666 14354
rect 1700 14320 1706 14354
rect 858 14306 1619 14312
rect 219 14272 231 14306
rect 1607 14272 1619 14306
rect 219 14266 352 14272
rect 132 14224 138 14258
rect 172 14224 178 14258
rect 342 14256 352 14266
rect 858 14266 1619 14272
rect 858 14256 868 14266
rect 132 14066 178 14224
rect 970 14216 980 14226
rect 219 14210 980 14216
rect 1490 14216 1500 14226
rect 1490 14210 1619 14216
rect 219 14176 231 14210
rect 1607 14176 1619 14210
rect 219 14170 980 14176
rect 970 14160 980 14170
rect 1490 14170 1619 14176
rect 1490 14160 1500 14170
rect 1660 14162 1706 14320
rect 342 14120 352 14130
rect 219 14114 352 14120
rect 858 14120 868 14130
rect 1660 14128 1666 14162
rect 1700 14128 1706 14162
rect 858 14114 1619 14120
rect 219 14080 231 14114
rect 1607 14080 1619 14114
rect 219 14074 352 14080
rect 132 14032 138 14066
rect 172 14032 178 14066
rect 342 14064 352 14074
rect 858 14074 1619 14080
rect 858 14064 868 14074
rect 132 13874 178 14032
rect 970 14024 980 14034
rect 219 14018 980 14024
rect 1490 14024 1500 14034
rect 1490 14018 1619 14024
rect 219 13984 231 14018
rect 1607 13984 1619 14018
rect 219 13978 980 13984
rect 970 13968 980 13978
rect 1490 13978 1619 13984
rect 1490 13968 1500 13978
rect 1660 13970 1706 14128
rect 342 13928 352 13938
rect 219 13922 352 13928
rect 858 13928 868 13938
rect 1660 13936 1666 13970
rect 1700 13936 1706 13970
rect 858 13922 1619 13928
rect 219 13888 231 13922
rect 1607 13888 1619 13922
rect 219 13882 352 13888
rect 132 13840 138 13874
rect 172 13840 178 13874
rect 342 13872 352 13882
rect 858 13882 1619 13888
rect 858 13872 868 13882
rect 132 13682 178 13840
rect 970 13832 980 13842
rect 219 13826 980 13832
rect 1490 13832 1500 13842
rect 1490 13826 1619 13832
rect 219 13792 231 13826
rect 1607 13792 1619 13826
rect 219 13786 980 13792
rect 970 13776 980 13786
rect 1490 13786 1619 13792
rect 1490 13776 1500 13786
rect 1660 13778 1706 13936
rect 342 13736 352 13746
rect 219 13730 352 13736
rect 858 13736 868 13746
rect 1660 13744 1666 13778
rect 1700 13744 1706 13778
rect 858 13730 1619 13736
rect 219 13696 231 13730
rect 1607 13696 1619 13730
rect 219 13690 352 13696
rect 132 13648 138 13682
rect 172 13648 178 13682
rect 342 13680 352 13690
rect 858 13690 1619 13696
rect 858 13680 868 13690
rect 132 13490 178 13648
rect 970 13640 980 13650
rect 219 13634 980 13640
rect 1490 13640 1500 13650
rect 1490 13634 1619 13640
rect 219 13600 231 13634
rect 1607 13600 1619 13634
rect 219 13594 980 13600
rect 970 13584 980 13594
rect 1490 13594 1619 13600
rect 1490 13584 1500 13594
rect 1660 13586 1706 13744
rect 342 13544 352 13554
rect 219 13538 352 13544
rect 858 13544 868 13554
rect 1660 13552 1666 13586
rect 1700 13552 1706 13586
rect 858 13538 1619 13544
rect 219 13504 231 13538
rect 1607 13504 1619 13538
rect 219 13498 352 13504
rect 132 13456 138 13490
rect 172 13456 178 13490
rect 342 13488 352 13498
rect 858 13498 1619 13504
rect 858 13488 868 13498
rect 132 13298 178 13456
rect 970 13448 980 13458
rect 219 13442 980 13448
rect 1490 13448 1500 13458
rect 1490 13442 1619 13448
rect 219 13408 231 13442
rect 1607 13408 1619 13442
rect 219 13402 980 13408
rect 970 13392 980 13402
rect 1490 13402 1619 13408
rect 1490 13392 1500 13402
rect 1660 13394 1706 13552
rect 342 13352 352 13362
rect 219 13346 352 13352
rect 858 13352 868 13362
rect 1660 13360 1666 13394
rect 1700 13360 1706 13394
rect 858 13346 1619 13352
rect 219 13312 231 13346
rect 1607 13312 1619 13346
rect 219 13306 352 13312
rect 132 13264 138 13298
rect 172 13264 178 13298
rect 342 13296 352 13306
rect 858 13306 1619 13312
rect 858 13296 868 13306
rect 132 13106 178 13264
rect 970 13256 980 13266
rect 219 13250 980 13256
rect 1490 13256 1500 13266
rect 1490 13250 1619 13256
rect 219 13216 231 13250
rect 1607 13216 1619 13250
rect 219 13210 980 13216
rect 970 13200 980 13210
rect 1490 13210 1619 13216
rect 1490 13200 1500 13210
rect 1660 13202 1706 13360
rect 342 13160 352 13170
rect 219 13154 352 13160
rect 858 13160 868 13170
rect 1660 13168 1666 13202
rect 1700 13168 1706 13202
rect 858 13154 1619 13160
rect 219 13120 231 13154
rect 1607 13120 1619 13154
rect 219 13114 352 13120
rect 132 13072 138 13106
rect 172 13072 178 13106
rect 342 13104 352 13114
rect 858 13114 1619 13120
rect 858 13104 868 13114
rect 132 12914 178 13072
rect 970 13064 980 13074
rect 219 13058 980 13064
rect 1490 13064 1500 13074
rect 1490 13058 1619 13064
rect 219 13024 231 13058
rect 1607 13024 1619 13058
rect 219 13018 980 13024
rect 970 13008 980 13018
rect 1490 13018 1619 13024
rect 1490 13008 1500 13018
rect 1660 13010 1706 13168
rect 342 12968 352 12978
rect 219 12962 352 12968
rect 858 12968 868 12978
rect 1660 12976 1666 13010
rect 1700 12976 1706 13010
rect 858 12962 1619 12968
rect 219 12928 231 12962
rect 1607 12928 1619 12962
rect 219 12922 352 12928
rect 132 12880 138 12914
rect 172 12880 178 12914
rect 342 12912 352 12922
rect 858 12922 1619 12928
rect 858 12912 868 12922
rect 132 12722 178 12880
rect 970 12872 980 12882
rect 219 12866 980 12872
rect 1490 12872 1500 12882
rect 1490 12866 1619 12872
rect 219 12832 231 12866
rect 1607 12832 1619 12866
rect 219 12826 980 12832
rect 970 12816 980 12826
rect 1490 12826 1619 12832
rect 1490 12816 1500 12826
rect 1660 12818 1706 12976
rect 342 12776 352 12786
rect 219 12770 352 12776
rect 858 12776 868 12786
rect 1660 12784 1666 12818
rect 1700 12784 1706 12818
rect 858 12770 1619 12776
rect 219 12736 231 12770
rect 1607 12736 1619 12770
rect 219 12730 352 12736
rect 132 12688 138 12722
rect 172 12688 178 12722
rect 342 12720 352 12730
rect 858 12730 1619 12736
rect 858 12720 868 12730
rect 132 12530 178 12688
rect 970 12680 980 12690
rect 219 12674 980 12680
rect 1490 12680 1500 12690
rect 1490 12674 1619 12680
rect 219 12640 231 12674
rect 1607 12640 1619 12674
rect 219 12634 980 12640
rect 970 12624 980 12634
rect 1490 12634 1619 12640
rect 1490 12624 1500 12634
rect 1660 12626 1706 12784
rect 342 12584 352 12594
rect 219 12578 352 12584
rect 858 12584 868 12594
rect 1660 12592 1666 12626
rect 1700 12592 1706 12626
rect 858 12578 1619 12584
rect 219 12544 231 12578
rect 1607 12544 1619 12578
rect 219 12538 352 12544
rect 132 12496 138 12530
rect 172 12496 178 12530
rect 342 12528 352 12538
rect 858 12538 1619 12544
rect 858 12528 868 12538
rect 132 12338 178 12496
rect 970 12488 980 12498
rect 219 12482 980 12488
rect 1490 12488 1500 12498
rect 1490 12482 1619 12488
rect 219 12448 231 12482
rect 1607 12448 1619 12482
rect 219 12442 980 12448
rect 970 12432 980 12442
rect 1490 12442 1619 12448
rect 1490 12432 1500 12442
rect 1660 12434 1706 12592
rect 342 12392 352 12402
rect 219 12386 352 12392
rect 858 12392 868 12402
rect 1660 12400 1666 12434
rect 1700 12400 1706 12434
rect 858 12386 1619 12392
rect 219 12352 231 12386
rect 1607 12352 1619 12386
rect 219 12346 352 12352
rect 132 12304 138 12338
rect 172 12304 178 12338
rect 342 12336 352 12346
rect 858 12346 1619 12352
rect 858 12336 868 12346
rect 132 12146 178 12304
rect 970 12296 980 12306
rect 219 12290 980 12296
rect 1490 12296 1500 12306
rect 1490 12290 1619 12296
rect 219 12256 231 12290
rect 1607 12256 1619 12290
rect 219 12250 980 12256
rect 970 12240 980 12250
rect 1490 12250 1619 12256
rect 1490 12240 1500 12250
rect 1660 12242 1706 12400
rect 342 12200 352 12210
rect 219 12194 352 12200
rect 858 12200 868 12210
rect 1660 12208 1666 12242
rect 1700 12208 1706 12242
rect 858 12194 1619 12200
rect 219 12160 231 12194
rect 1607 12160 1619 12194
rect 219 12154 352 12160
rect 132 12112 138 12146
rect 172 12112 178 12146
rect 342 12144 352 12154
rect 858 12154 1619 12160
rect 858 12144 868 12154
rect 132 11954 178 12112
rect 970 12104 980 12114
rect 219 12098 980 12104
rect 1490 12104 1500 12114
rect 1490 12098 1619 12104
rect 219 12064 231 12098
rect 1607 12064 1619 12098
rect 219 12058 980 12064
rect 970 12048 980 12058
rect 1490 12058 1619 12064
rect 1490 12048 1500 12058
rect 1660 12050 1706 12208
rect 342 12008 352 12018
rect 219 12002 352 12008
rect 858 12008 868 12018
rect 1660 12016 1666 12050
rect 1700 12016 1706 12050
rect 858 12002 1619 12008
rect 219 11968 231 12002
rect 1607 11968 1619 12002
rect 219 11962 352 11968
rect 132 11920 138 11954
rect 172 11920 178 11954
rect 342 11952 352 11962
rect 858 11962 1619 11968
rect 858 11952 868 11962
rect 132 11762 178 11920
rect 970 11912 980 11922
rect 219 11906 980 11912
rect 1490 11912 1500 11922
rect 1490 11906 1619 11912
rect 219 11872 231 11906
rect 1607 11872 1619 11906
rect 219 11866 980 11872
rect 970 11856 980 11866
rect 1490 11866 1619 11872
rect 1490 11856 1500 11866
rect 1660 11858 1706 12016
rect 342 11816 352 11826
rect 219 11810 352 11816
rect 858 11816 868 11826
rect 1660 11824 1666 11858
rect 1700 11824 1706 11858
rect 858 11810 1619 11816
rect 219 11776 231 11810
rect 1607 11776 1619 11810
rect 219 11770 352 11776
rect 132 11728 138 11762
rect 172 11728 178 11762
rect 342 11760 352 11770
rect 858 11770 1619 11776
rect 858 11760 868 11770
rect 132 11570 178 11728
rect 970 11720 980 11730
rect 219 11714 980 11720
rect 1490 11720 1500 11730
rect 1490 11714 1619 11720
rect 219 11680 231 11714
rect 1607 11680 1619 11714
rect 219 11674 980 11680
rect 970 11664 980 11674
rect 1490 11674 1619 11680
rect 1490 11664 1500 11674
rect 1660 11666 1706 11824
rect 342 11624 352 11634
rect 219 11618 352 11624
rect 858 11624 868 11634
rect 1660 11632 1666 11666
rect 1700 11632 1706 11666
rect 858 11618 1619 11624
rect 219 11584 231 11618
rect 1607 11584 1619 11618
rect 219 11578 352 11584
rect 132 11536 138 11570
rect 172 11536 178 11570
rect 342 11568 352 11578
rect 858 11578 1619 11584
rect 858 11568 868 11578
rect 132 11378 178 11536
rect 970 11528 980 11538
rect 219 11522 980 11528
rect 1490 11528 1500 11538
rect 1490 11522 1619 11528
rect 219 11488 231 11522
rect 1607 11488 1619 11522
rect 219 11482 980 11488
rect 970 11472 980 11482
rect 1490 11482 1619 11488
rect 1490 11472 1500 11482
rect 1660 11474 1706 11632
rect 342 11432 352 11442
rect 219 11426 352 11432
rect 858 11432 868 11442
rect 1660 11440 1666 11474
rect 1700 11440 1706 11474
rect 858 11426 1619 11432
rect 219 11392 231 11426
rect 1607 11392 1619 11426
rect 219 11386 352 11392
rect 132 11344 138 11378
rect 172 11344 178 11378
rect 342 11376 352 11386
rect 858 11386 1619 11392
rect 858 11376 868 11386
rect 132 11186 178 11344
rect 970 11336 980 11346
rect 219 11330 980 11336
rect 1490 11336 1500 11346
rect 1490 11330 1619 11336
rect 219 11296 231 11330
rect 1607 11296 1619 11330
rect 219 11290 980 11296
rect 970 11280 980 11290
rect 1490 11290 1619 11296
rect 1490 11280 1500 11290
rect 1660 11282 1706 11440
rect 342 11240 352 11250
rect 219 11234 352 11240
rect 858 11240 868 11250
rect 1660 11248 1666 11282
rect 1700 11248 1706 11282
rect 858 11234 1619 11240
rect 219 11200 231 11234
rect 1607 11200 1619 11234
rect 219 11194 352 11200
rect 132 11152 138 11186
rect 172 11152 178 11186
rect 342 11184 352 11194
rect 858 11194 1619 11200
rect 858 11184 868 11194
rect 132 10994 178 11152
rect 970 11144 980 11154
rect 219 11138 980 11144
rect 1490 11144 1500 11154
rect 1490 11138 1619 11144
rect 219 11104 231 11138
rect 1607 11104 1619 11138
rect 219 11098 980 11104
rect 970 11088 980 11098
rect 1490 11098 1619 11104
rect 1490 11088 1500 11098
rect 1660 11090 1706 11248
rect 342 11048 352 11058
rect 219 11042 352 11048
rect 858 11048 868 11058
rect 1660 11056 1666 11090
rect 1700 11056 1706 11090
rect 858 11042 1619 11048
rect 219 11008 231 11042
rect 1607 11008 1619 11042
rect 219 11002 352 11008
rect 132 10960 138 10994
rect 172 10960 178 10994
rect 342 10992 352 11002
rect 858 11002 1619 11008
rect 858 10992 868 11002
rect 132 10802 178 10960
rect 970 10952 980 10962
rect 219 10946 980 10952
rect 1490 10952 1500 10962
rect 1490 10946 1619 10952
rect 219 10912 231 10946
rect 1607 10912 1619 10946
rect 219 10906 980 10912
rect 970 10896 980 10906
rect 1490 10906 1619 10912
rect 1490 10896 1500 10906
rect 1660 10898 1706 11056
rect 342 10856 352 10866
rect 219 10850 352 10856
rect 858 10856 868 10866
rect 1660 10864 1666 10898
rect 1700 10864 1706 10898
rect 858 10850 1619 10856
rect 219 10816 231 10850
rect 1607 10816 1619 10850
rect 219 10810 352 10816
rect 132 10768 138 10802
rect 172 10768 178 10802
rect 342 10800 352 10810
rect 858 10810 1619 10816
rect 858 10800 868 10810
rect 132 10610 178 10768
rect 970 10760 980 10770
rect 219 10754 980 10760
rect 1490 10760 1500 10770
rect 1490 10754 1619 10760
rect 219 10720 231 10754
rect 1607 10720 1619 10754
rect 219 10714 980 10720
rect 970 10704 980 10714
rect 1490 10714 1619 10720
rect 1490 10704 1500 10714
rect 1660 10706 1706 10864
rect 342 10664 352 10674
rect 219 10658 352 10664
rect 858 10664 868 10674
rect 1660 10672 1666 10706
rect 1700 10672 1706 10706
rect 858 10658 1619 10664
rect 219 10624 231 10658
rect 1607 10624 1619 10658
rect 219 10618 352 10624
rect 132 10576 138 10610
rect 172 10576 178 10610
rect 342 10608 352 10618
rect 858 10618 1619 10624
rect 858 10608 868 10618
rect 132 10418 178 10576
rect 970 10568 980 10578
rect 219 10562 980 10568
rect 1490 10568 1500 10578
rect 1490 10562 1619 10568
rect 219 10528 231 10562
rect 1607 10528 1619 10562
rect 219 10522 980 10528
rect 970 10512 980 10522
rect 1490 10522 1619 10528
rect 1490 10512 1500 10522
rect 1660 10514 1706 10672
rect 342 10472 352 10482
rect 219 10466 352 10472
rect 858 10472 868 10482
rect 1660 10480 1666 10514
rect 1700 10480 1706 10514
rect 858 10466 1619 10472
rect 219 10432 231 10466
rect 1607 10432 1619 10466
rect 219 10426 352 10432
rect 132 10384 138 10418
rect 172 10384 178 10418
rect 342 10416 352 10426
rect 858 10426 1619 10432
rect 858 10416 868 10426
rect 132 10226 178 10384
rect 970 10376 980 10386
rect 219 10370 980 10376
rect 1490 10376 1500 10386
rect 1490 10370 1619 10376
rect 219 10336 231 10370
rect 1607 10336 1619 10370
rect 219 10330 980 10336
rect 970 10320 980 10330
rect 1490 10330 1619 10336
rect 1490 10320 1500 10330
rect 1660 10322 1706 10480
rect 342 10280 352 10290
rect 219 10274 352 10280
rect 858 10280 868 10290
rect 1660 10288 1666 10322
rect 1700 10288 1706 10322
rect 858 10274 1619 10280
rect 219 10240 231 10274
rect 1607 10240 1619 10274
rect 219 10234 352 10240
rect 132 10192 138 10226
rect 172 10192 178 10226
rect 342 10224 352 10234
rect 858 10234 1619 10240
rect 858 10224 868 10234
rect 132 10034 178 10192
rect 970 10184 980 10194
rect 219 10178 980 10184
rect 1490 10184 1500 10194
rect 1490 10178 1619 10184
rect 219 10144 231 10178
rect 1607 10144 1619 10178
rect 219 10138 980 10144
rect 970 10128 980 10138
rect 1490 10138 1619 10144
rect 1490 10128 1500 10138
rect 1660 10130 1706 10288
rect 342 10088 352 10098
rect 219 10082 352 10088
rect 858 10088 868 10098
rect 1660 10096 1666 10130
rect 1700 10096 1706 10130
rect 858 10082 1619 10088
rect 219 10048 231 10082
rect 1607 10048 1619 10082
rect 219 10042 352 10048
rect 132 10000 138 10034
rect 172 10000 178 10034
rect 342 10032 352 10042
rect 858 10042 1619 10048
rect 858 10032 868 10042
rect 132 9842 178 10000
rect 970 9992 980 10002
rect 219 9986 980 9992
rect 1490 9992 1500 10002
rect 1490 9986 1619 9992
rect 219 9952 231 9986
rect 1607 9952 1619 9986
rect 219 9946 980 9952
rect 970 9936 980 9946
rect 1490 9946 1619 9952
rect 1490 9936 1500 9946
rect 1660 9938 1706 10096
rect 342 9896 352 9906
rect 219 9890 352 9896
rect 858 9896 868 9906
rect 1660 9904 1666 9938
rect 1700 9904 1706 9938
rect 858 9890 1619 9896
rect 219 9856 231 9890
rect 1607 9856 1619 9890
rect 219 9850 352 9856
rect 132 9808 138 9842
rect 172 9808 178 9842
rect 342 9840 352 9850
rect 858 9850 1619 9856
rect 858 9840 868 9850
rect 132 9650 178 9808
rect 970 9800 980 9810
rect 219 9794 980 9800
rect 1490 9800 1500 9810
rect 1490 9794 1619 9800
rect 219 9760 231 9794
rect 1607 9760 1619 9794
rect 219 9754 980 9760
rect 970 9744 980 9754
rect 1490 9754 1619 9760
rect 1490 9744 1500 9754
rect 1660 9746 1706 9904
rect 342 9704 352 9714
rect 219 9698 352 9704
rect 858 9704 868 9714
rect 1660 9712 1666 9746
rect 1700 9712 1706 9746
rect 858 9698 1619 9704
rect 219 9664 231 9698
rect 1607 9664 1619 9698
rect 219 9658 352 9664
rect 132 9616 138 9650
rect 172 9616 178 9650
rect 342 9648 352 9658
rect 858 9658 1619 9664
rect 858 9648 868 9658
rect 132 9458 178 9616
rect 970 9608 980 9618
rect 219 9602 980 9608
rect 1490 9608 1500 9618
rect 1490 9602 1619 9608
rect 219 9568 231 9602
rect 1607 9568 1619 9602
rect 219 9562 980 9568
rect 970 9552 980 9562
rect 1490 9562 1619 9568
rect 1490 9552 1500 9562
rect 1660 9554 1706 9712
rect 342 9512 352 9522
rect 219 9506 352 9512
rect 858 9512 868 9522
rect 1660 9520 1666 9554
rect 1700 9520 1706 9554
rect 858 9506 1619 9512
rect 219 9472 231 9506
rect 1607 9472 1619 9506
rect 219 9466 352 9472
rect 132 9424 138 9458
rect 172 9424 178 9458
rect 342 9456 352 9466
rect 858 9466 1619 9472
rect 858 9456 868 9466
rect 132 9266 178 9424
rect 970 9416 980 9426
rect 219 9410 980 9416
rect 1490 9416 1500 9426
rect 1490 9410 1619 9416
rect 219 9376 231 9410
rect 1607 9376 1619 9410
rect 219 9370 980 9376
rect 970 9360 980 9370
rect 1490 9370 1619 9376
rect 1490 9360 1500 9370
rect 1660 9362 1706 9520
rect 342 9320 352 9330
rect 219 9314 352 9320
rect 858 9320 868 9330
rect 1660 9328 1666 9362
rect 1700 9328 1706 9362
rect 858 9314 1619 9320
rect 219 9280 231 9314
rect 1607 9280 1619 9314
rect 219 9274 352 9280
rect 132 9232 138 9266
rect 172 9232 178 9266
rect 342 9264 352 9274
rect 858 9274 1619 9280
rect 858 9264 868 9274
rect 132 9074 178 9232
rect 970 9224 980 9234
rect 219 9218 980 9224
rect 1490 9224 1500 9234
rect 1490 9218 1619 9224
rect 219 9184 231 9218
rect 1607 9184 1619 9218
rect 219 9178 980 9184
rect 970 9168 980 9178
rect 1490 9178 1619 9184
rect 1490 9168 1500 9178
rect 1660 9170 1706 9328
rect 342 9128 352 9138
rect 219 9122 352 9128
rect 858 9128 868 9138
rect 1660 9136 1666 9170
rect 1700 9136 1706 9170
rect 858 9122 1619 9128
rect 219 9088 231 9122
rect 1607 9088 1619 9122
rect 219 9082 352 9088
rect 132 9040 138 9074
rect 172 9040 178 9074
rect 342 9072 352 9082
rect 858 9082 1619 9088
rect 858 9072 868 9082
rect 132 8882 178 9040
rect 970 9032 980 9042
rect 219 9026 980 9032
rect 1490 9032 1500 9042
rect 1490 9026 1619 9032
rect 219 8992 231 9026
rect 1607 8992 1619 9026
rect 219 8986 980 8992
rect 970 8976 980 8986
rect 1490 8986 1619 8992
rect 1490 8976 1500 8986
rect 1660 8978 1706 9136
rect 342 8936 352 8946
rect 219 8930 352 8936
rect 858 8936 868 8946
rect 1660 8944 1666 8978
rect 1700 8944 1706 8978
rect 858 8930 1619 8936
rect 219 8896 231 8930
rect 1607 8896 1619 8930
rect 219 8890 352 8896
rect 132 8848 138 8882
rect 172 8848 178 8882
rect 342 8880 352 8890
rect 858 8890 1619 8896
rect 858 8880 868 8890
rect 132 8690 178 8848
rect 970 8840 980 8850
rect 219 8834 980 8840
rect 1490 8840 1500 8850
rect 1490 8834 1619 8840
rect 219 8800 231 8834
rect 1607 8800 1619 8834
rect 219 8794 980 8800
rect 970 8784 980 8794
rect 1490 8794 1619 8800
rect 1490 8784 1500 8794
rect 1660 8786 1706 8944
rect 342 8744 352 8754
rect 219 8738 352 8744
rect 858 8744 868 8754
rect 1660 8752 1666 8786
rect 1700 8752 1706 8786
rect 858 8738 1619 8744
rect 219 8704 231 8738
rect 1607 8704 1619 8738
rect 219 8698 352 8704
rect 132 8656 138 8690
rect 172 8656 178 8690
rect 342 8688 352 8698
rect 858 8698 1619 8704
rect 858 8688 868 8698
rect 132 8498 178 8656
rect 970 8648 980 8658
rect 219 8642 980 8648
rect 1490 8648 1500 8658
rect 1490 8642 1619 8648
rect 219 8608 231 8642
rect 1607 8608 1619 8642
rect 219 8602 980 8608
rect 970 8592 980 8602
rect 1490 8602 1619 8608
rect 1490 8592 1500 8602
rect 1660 8594 1706 8752
rect 342 8552 352 8562
rect 219 8546 352 8552
rect 858 8552 868 8562
rect 1660 8560 1666 8594
rect 1700 8560 1706 8594
rect 858 8546 1619 8552
rect 219 8512 231 8546
rect 1607 8512 1619 8546
rect 219 8506 352 8512
rect 132 8464 138 8498
rect 172 8464 178 8498
rect 342 8496 352 8506
rect 858 8506 1619 8512
rect 858 8496 868 8506
rect 132 8306 178 8464
rect 970 8456 980 8466
rect 219 8450 980 8456
rect 1490 8456 1500 8466
rect 1490 8450 1619 8456
rect 219 8416 231 8450
rect 1607 8416 1619 8450
rect 219 8410 980 8416
rect 970 8400 980 8410
rect 1490 8410 1619 8416
rect 1490 8400 1500 8410
rect 1660 8402 1706 8560
rect 342 8360 352 8370
rect 219 8354 352 8360
rect 858 8360 868 8370
rect 1660 8368 1666 8402
rect 1700 8368 1706 8402
rect 858 8354 1619 8360
rect 219 8320 231 8354
rect 1607 8320 1619 8354
rect 219 8314 352 8320
rect 132 8272 138 8306
rect 172 8272 178 8306
rect 342 8304 352 8314
rect 858 8314 1619 8320
rect 858 8304 868 8314
rect 132 8114 178 8272
rect 970 8264 980 8274
rect 219 8258 980 8264
rect 1490 8264 1500 8274
rect 1490 8258 1619 8264
rect 219 8224 231 8258
rect 1607 8224 1619 8258
rect 219 8218 980 8224
rect 970 8208 980 8218
rect 1490 8218 1619 8224
rect 1490 8208 1500 8218
rect 1660 8210 1706 8368
rect 342 8168 352 8178
rect 219 8162 352 8168
rect 858 8168 868 8178
rect 1660 8176 1666 8210
rect 1700 8176 1706 8210
rect 858 8162 1619 8168
rect 219 8128 231 8162
rect 1607 8128 1619 8162
rect 219 8122 352 8128
rect 132 8080 138 8114
rect 172 8080 178 8114
rect 342 8112 352 8122
rect 858 8122 1619 8128
rect 858 8112 868 8122
rect 132 7922 178 8080
rect 970 8072 980 8082
rect 219 8066 980 8072
rect 1490 8072 1500 8082
rect 1490 8066 1619 8072
rect 219 8032 231 8066
rect 1607 8032 1619 8066
rect 219 8026 980 8032
rect 970 8016 980 8026
rect 1490 8026 1619 8032
rect 1490 8016 1500 8026
rect 1660 8018 1706 8176
rect 342 7976 352 7986
rect 219 7970 352 7976
rect 858 7976 868 7986
rect 1660 7984 1666 8018
rect 1700 7984 1706 8018
rect 858 7970 1619 7976
rect 219 7936 231 7970
rect 1607 7936 1619 7970
rect 219 7930 352 7936
rect 132 7888 138 7922
rect 172 7888 178 7922
rect 342 7920 352 7930
rect 858 7930 1619 7936
rect 858 7920 868 7930
rect 132 7730 178 7888
rect 970 7880 980 7890
rect 219 7874 980 7880
rect 1490 7880 1500 7890
rect 1490 7874 1619 7880
rect 219 7840 231 7874
rect 1607 7840 1619 7874
rect 219 7834 980 7840
rect 970 7824 980 7834
rect 1490 7834 1619 7840
rect 1490 7824 1500 7834
rect 1660 7826 1706 7984
rect 342 7784 352 7794
rect 219 7778 352 7784
rect 858 7784 868 7794
rect 1660 7792 1666 7826
rect 1700 7792 1706 7826
rect 858 7778 1619 7784
rect 219 7744 231 7778
rect 1607 7744 1619 7778
rect 219 7738 352 7744
rect 132 7696 138 7730
rect 172 7696 178 7730
rect 342 7728 352 7738
rect 858 7738 1619 7744
rect 858 7728 868 7738
rect 132 7538 178 7696
rect 970 7688 980 7698
rect 219 7682 980 7688
rect 1490 7688 1500 7698
rect 1490 7682 1619 7688
rect 219 7648 231 7682
rect 1607 7648 1619 7682
rect 219 7642 980 7648
rect 970 7632 980 7642
rect 1490 7642 1619 7648
rect 1490 7632 1500 7642
rect 1660 7634 1706 7792
rect 342 7592 352 7602
rect 219 7586 352 7592
rect 858 7592 868 7602
rect 1660 7600 1666 7634
rect 1700 7600 1706 7634
rect 858 7586 1619 7592
rect 219 7552 231 7586
rect 1607 7552 1619 7586
rect 219 7546 352 7552
rect 132 7504 138 7538
rect 172 7504 178 7538
rect 342 7536 352 7546
rect 858 7546 1619 7552
rect 858 7536 868 7546
rect 132 7346 178 7504
rect 970 7496 980 7506
rect 219 7490 980 7496
rect 1490 7496 1500 7506
rect 1490 7490 1619 7496
rect 219 7456 231 7490
rect 1607 7456 1619 7490
rect 219 7450 980 7456
rect 970 7440 980 7450
rect 1490 7450 1619 7456
rect 1490 7440 1500 7450
rect 1660 7442 1706 7600
rect 342 7400 352 7410
rect 219 7394 352 7400
rect 858 7400 868 7410
rect 1660 7408 1666 7442
rect 1700 7408 1706 7442
rect 858 7394 1619 7400
rect 219 7360 231 7394
rect 1607 7360 1619 7394
rect 219 7354 352 7360
rect 132 7312 138 7346
rect 172 7312 178 7346
rect 342 7344 352 7354
rect 858 7354 1619 7360
rect 858 7344 868 7354
rect 132 7154 178 7312
rect 970 7304 980 7314
rect 219 7298 980 7304
rect 1490 7304 1500 7314
rect 1490 7298 1619 7304
rect 219 7264 231 7298
rect 1607 7264 1619 7298
rect 219 7258 980 7264
rect 970 7248 980 7258
rect 1490 7258 1619 7264
rect 1490 7248 1500 7258
rect 1660 7250 1706 7408
rect 342 7208 352 7218
rect 219 7202 352 7208
rect 858 7208 868 7218
rect 1660 7216 1666 7250
rect 1700 7216 1706 7250
rect 858 7202 1619 7208
rect 219 7168 231 7202
rect 1607 7168 1619 7202
rect 219 7162 352 7168
rect 132 7120 138 7154
rect 172 7120 178 7154
rect 342 7152 352 7162
rect 858 7162 1619 7168
rect 858 7152 868 7162
rect 132 6962 178 7120
rect 970 7112 980 7122
rect 219 7106 980 7112
rect 1490 7112 1500 7122
rect 1490 7106 1619 7112
rect 219 7072 231 7106
rect 1607 7072 1619 7106
rect 219 7066 980 7072
rect 970 7056 980 7066
rect 1490 7066 1619 7072
rect 1490 7056 1500 7066
rect 1660 7058 1706 7216
rect 342 7016 352 7026
rect 219 7010 352 7016
rect 858 7016 868 7026
rect 1660 7024 1666 7058
rect 1700 7024 1706 7058
rect 858 7010 1619 7016
rect 219 6976 231 7010
rect 1607 6976 1619 7010
rect 219 6970 352 6976
rect 132 6928 138 6962
rect 172 6928 178 6962
rect 342 6960 352 6970
rect 858 6970 1619 6976
rect 858 6960 868 6970
rect 132 6770 178 6928
rect 970 6920 980 6930
rect 219 6914 980 6920
rect 1490 6920 1500 6930
rect 1490 6914 1619 6920
rect 219 6880 231 6914
rect 1607 6880 1619 6914
rect 219 6874 980 6880
rect 970 6864 980 6874
rect 1490 6874 1619 6880
rect 1490 6864 1500 6874
rect 1660 6866 1706 7024
rect 342 6824 352 6834
rect 219 6818 352 6824
rect 858 6824 868 6834
rect 1660 6832 1666 6866
rect 1700 6832 1706 6866
rect 858 6818 1619 6824
rect 219 6784 231 6818
rect 1607 6784 1619 6818
rect 219 6778 352 6784
rect 132 6736 138 6770
rect 172 6736 178 6770
rect 342 6768 352 6778
rect 858 6778 1619 6784
rect 858 6768 868 6778
rect 132 6578 178 6736
rect 970 6728 980 6738
rect 219 6722 980 6728
rect 1490 6728 1500 6738
rect 1490 6722 1619 6728
rect 219 6688 231 6722
rect 1607 6688 1619 6722
rect 219 6682 980 6688
rect 970 6672 980 6682
rect 1490 6682 1619 6688
rect 1490 6672 1500 6682
rect 1660 6674 1706 6832
rect 342 6632 352 6642
rect 219 6626 352 6632
rect 858 6632 868 6642
rect 1660 6640 1666 6674
rect 1700 6640 1706 6674
rect 858 6626 1619 6632
rect 219 6592 231 6626
rect 1607 6592 1619 6626
rect 219 6586 352 6592
rect 132 6544 138 6578
rect 172 6544 178 6578
rect 342 6576 352 6586
rect 858 6586 1619 6592
rect 858 6576 868 6586
rect 132 6386 178 6544
rect 970 6536 980 6546
rect 219 6530 980 6536
rect 1490 6536 1500 6546
rect 1490 6530 1619 6536
rect 219 6496 231 6530
rect 1607 6496 1619 6530
rect 219 6490 980 6496
rect 970 6480 980 6490
rect 1490 6490 1619 6496
rect 1490 6480 1500 6490
rect 1660 6482 1706 6640
rect 342 6440 352 6450
rect 219 6434 352 6440
rect 858 6440 868 6450
rect 1660 6448 1666 6482
rect 1700 6448 1706 6482
rect 858 6434 1619 6440
rect 219 6400 231 6434
rect 1607 6400 1619 6434
rect 219 6394 352 6400
rect 132 6352 138 6386
rect 172 6352 178 6386
rect 342 6384 352 6394
rect 858 6394 1619 6400
rect 858 6384 868 6394
rect 132 6194 178 6352
rect 970 6344 980 6354
rect 219 6338 980 6344
rect 1490 6344 1500 6354
rect 1490 6338 1619 6344
rect 219 6304 231 6338
rect 1607 6304 1619 6338
rect 219 6298 980 6304
rect 970 6288 980 6298
rect 1490 6298 1619 6304
rect 1490 6288 1500 6298
rect 1660 6290 1706 6448
rect 342 6248 352 6258
rect 219 6242 352 6248
rect 858 6248 868 6258
rect 1660 6256 1666 6290
rect 1700 6256 1706 6290
rect 858 6242 1619 6248
rect 219 6208 231 6242
rect 1607 6208 1619 6242
rect 219 6202 352 6208
rect 132 6160 138 6194
rect 172 6160 178 6194
rect 342 6192 352 6202
rect 858 6202 1619 6208
rect 858 6192 868 6202
rect 132 6002 178 6160
rect 970 6152 980 6162
rect 219 6146 980 6152
rect 1490 6152 1500 6162
rect 1490 6146 1619 6152
rect 219 6112 231 6146
rect 1607 6112 1619 6146
rect 219 6106 980 6112
rect 970 6096 980 6106
rect 1490 6106 1619 6112
rect 1490 6096 1500 6106
rect 1660 6098 1706 6256
rect 342 6056 352 6066
rect 219 6050 352 6056
rect 858 6056 868 6066
rect 1660 6064 1666 6098
rect 1700 6064 1706 6098
rect 858 6050 1619 6056
rect 219 6016 231 6050
rect 1607 6016 1619 6050
rect 219 6010 352 6016
rect 132 5968 138 6002
rect 172 5968 178 6002
rect 342 6000 352 6010
rect 858 6010 1619 6016
rect 858 6000 868 6010
rect 132 5810 178 5968
rect 970 5960 980 5970
rect 219 5954 980 5960
rect 1490 5960 1500 5970
rect 1490 5954 1619 5960
rect 219 5920 231 5954
rect 1607 5920 1619 5954
rect 219 5914 980 5920
rect 970 5904 980 5914
rect 1490 5914 1619 5920
rect 1490 5904 1500 5914
rect 1660 5906 1706 6064
rect 342 5864 352 5874
rect 219 5858 352 5864
rect 858 5864 868 5874
rect 1660 5872 1666 5906
rect 1700 5872 1706 5906
rect 858 5858 1619 5864
rect 219 5824 231 5858
rect 1607 5824 1619 5858
rect 219 5818 352 5824
rect 132 5776 138 5810
rect 172 5776 178 5810
rect 342 5808 352 5818
rect 858 5818 1619 5824
rect 858 5808 868 5818
rect 132 5618 178 5776
rect 970 5768 980 5778
rect 219 5762 980 5768
rect 1490 5768 1500 5778
rect 1490 5762 1619 5768
rect 219 5728 231 5762
rect 1607 5728 1619 5762
rect 219 5722 980 5728
rect 970 5712 980 5722
rect 1490 5722 1619 5728
rect 1490 5712 1500 5722
rect 1660 5714 1706 5872
rect 342 5672 352 5682
rect 219 5666 352 5672
rect 858 5672 868 5682
rect 1660 5680 1666 5714
rect 1700 5680 1706 5714
rect 858 5666 1619 5672
rect 219 5632 231 5666
rect 1607 5632 1619 5666
rect 219 5626 352 5632
rect 132 5584 138 5618
rect 172 5584 178 5618
rect 342 5616 352 5626
rect 858 5626 1619 5632
rect 858 5616 868 5626
rect 132 5426 178 5584
rect 970 5576 980 5586
rect 219 5570 980 5576
rect 1490 5576 1500 5586
rect 1490 5570 1619 5576
rect 219 5536 231 5570
rect 1607 5536 1619 5570
rect 219 5530 980 5536
rect 970 5520 980 5530
rect 1490 5530 1619 5536
rect 1490 5520 1500 5530
rect 1660 5522 1706 5680
rect 342 5480 352 5490
rect 219 5474 352 5480
rect 858 5480 868 5490
rect 1660 5488 1666 5522
rect 1700 5488 1706 5522
rect 858 5474 1619 5480
rect 219 5440 231 5474
rect 1607 5440 1619 5474
rect 219 5434 352 5440
rect 132 5392 138 5426
rect 172 5392 178 5426
rect 342 5424 352 5434
rect 858 5434 1619 5440
rect 858 5424 868 5434
rect 132 5234 178 5392
rect 970 5384 980 5394
rect 219 5378 980 5384
rect 1490 5384 1500 5394
rect 1490 5378 1619 5384
rect 219 5344 231 5378
rect 1607 5344 1619 5378
rect 219 5338 980 5344
rect 970 5328 980 5338
rect 1490 5338 1619 5344
rect 1490 5328 1500 5338
rect 1660 5330 1706 5488
rect 342 5288 352 5298
rect 219 5282 352 5288
rect 858 5288 868 5298
rect 1660 5296 1666 5330
rect 1700 5296 1706 5330
rect 858 5282 1619 5288
rect 219 5248 231 5282
rect 1607 5248 1619 5282
rect 219 5242 352 5248
rect 132 5200 138 5234
rect 172 5200 178 5234
rect 342 5232 352 5242
rect 858 5242 1619 5248
rect 858 5232 868 5242
rect 132 5042 178 5200
rect 970 5192 980 5202
rect 219 5186 980 5192
rect 1490 5192 1500 5202
rect 1490 5186 1619 5192
rect 219 5152 231 5186
rect 1607 5152 1619 5186
rect 219 5146 980 5152
rect 970 5136 980 5146
rect 1490 5146 1619 5152
rect 1490 5136 1500 5146
rect 1660 5138 1706 5296
rect 342 5096 352 5106
rect 219 5090 352 5096
rect 858 5096 868 5106
rect 1660 5104 1666 5138
rect 1700 5104 1706 5138
rect 858 5090 1619 5096
rect 219 5056 231 5090
rect 1607 5056 1619 5090
rect 219 5050 352 5056
rect 132 5008 138 5042
rect 172 5008 178 5042
rect 342 5040 352 5050
rect 858 5050 1619 5056
rect 858 5040 868 5050
rect 132 4850 178 5008
rect 970 5000 980 5010
rect 219 4994 980 5000
rect 1490 5000 1500 5010
rect 1490 4994 1619 5000
rect 219 4960 231 4994
rect 1607 4960 1619 4994
rect 219 4954 980 4960
rect 970 4944 980 4954
rect 1490 4954 1619 4960
rect 1490 4944 1500 4954
rect 1660 4946 1706 5104
rect 342 4904 352 4914
rect 219 4898 352 4904
rect 858 4904 868 4914
rect 1660 4912 1666 4946
rect 1700 4912 1706 4946
rect 858 4898 1619 4904
rect 219 4864 231 4898
rect 1607 4864 1619 4898
rect 219 4858 352 4864
rect 132 4816 138 4850
rect 172 4816 178 4850
rect 342 4848 352 4858
rect 858 4858 1619 4864
rect 858 4848 868 4858
rect 132 4658 178 4816
rect 970 4808 980 4818
rect 219 4802 980 4808
rect 1490 4808 1500 4818
rect 1490 4802 1619 4808
rect 219 4768 231 4802
rect 1607 4768 1619 4802
rect 219 4762 980 4768
rect 970 4752 980 4762
rect 1490 4762 1619 4768
rect 1490 4752 1500 4762
rect 1660 4754 1706 4912
rect 342 4712 352 4722
rect 219 4706 352 4712
rect 858 4712 868 4722
rect 1660 4720 1666 4754
rect 1700 4720 1706 4754
rect 858 4706 1619 4712
rect 219 4672 231 4706
rect 1607 4672 1619 4706
rect 219 4666 352 4672
rect 132 4624 138 4658
rect 172 4624 178 4658
rect 342 4656 352 4666
rect 858 4666 1619 4672
rect 858 4656 868 4666
rect 132 4466 178 4624
rect 970 4616 980 4626
rect 219 4610 980 4616
rect 1490 4616 1500 4626
rect 1490 4610 1619 4616
rect 219 4576 231 4610
rect 1607 4576 1619 4610
rect 219 4570 980 4576
rect 970 4560 980 4570
rect 1490 4570 1619 4576
rect 1490 4560 1500 4570
rect 1660 4562 1706 4720
rect 342 4520 352 4530
rect 219 4514 352 4520
rect 858 4520 868 4530
rect 1660 4528 1666 4562
rect 1700 4528 1706 4562
rect 858 4514 1619 4520
rect 219 4480 231 4514
rect 1607 4480 1619 4514
rect 219 4474 352 4480
rect 132 4432 138 4466
rect 172 4432 178 4466
rect 342 4464 352 4474
rect 858 4474 1619 4480
rect 858 4464 868 4474
rect 132 4274 178 4432
rect 970 4424 980 4434
rect 219 4418 980 4424
rect 1490 4424 1500 4434
rect 1490 4418 1619 4424
rect 219 4384 231 4418
rect 1607 4384 1619 4418
rect 219 4378 980 4384
rect 970 4368 980 4378
rect 1490 4378 1619 4384
rect 1490 4368 1500 4378
rect 1660 4370 1706 4528
rect 342 4328 352 4338
rect 219 4322 352 4328
rect 858 4328 868 4338
rect 1660 4336 1666 4370
rect 1700 4336 1706 4370
rect 858 4322 1619 4328
rect 219 4288 231 4322
rect 1607 4288 1619 4322
rect 219 4282 352 4288
rect 132 4240 138 4274
rect 172 4240 178 4274
rect 342 4272 352 4282
rect 858 4282 1619 4288
rect 858 4272 868 4282
rect 132 4082 178 4240
rect 970 4232 980 4242
rect 219 4226 980 4232
rect 1490 4232 1500 4242
rect 1490 4226 1619 4232
rect 219 4192 231 4226
rect 1607 4192 1619 4226
rect 219 4186 980 4192
rect 970 4176 980 4186
rect 1490 4186 1619 4192
rect 1490 4176 1500 4186
rect 1660 4178 1706 4336
rect 342 4136 352 4146
rect 219 4130 352 4136
rect 858 4136 868 4146
rect 1660 4144 1666 4178
rect 1700 4144 1706 4178
rect 858 4130 1619 4136
rect 219 4096 231 4130
rect 1607 4096 1619 4130
rect 219 4090 352 4096
rect 132 4048 138 4082
rect 172 4048 178 4082
rect 342 4080 352 4090
rect 858 4090 1619 4096
rect 858 4080 868 4090
rect 132 3890 178 4048
rect 970 4040 980 4050
rect 219 4034 980 4040
rect 1490 4040 1500 4050
rect 1490 4034 1619 4040
rect 219 4000 231 4034
rect 1607 4000 1619 4034
rect 219 3994 980 4000
rect 970 3984 980 3994
rect 1490 3994 1619 4000
rect 1490 3984 1500 3994
rect 1660 3986 1706 4144
rect 342 3944 352 3954
rect 219 3938 352 3944
rect 858 3944 868 3954
rect 1660 3952 1666 3986
rect 1700 3952 1706 3986
rect 858 3938 1619 3944
rect 219 3904 231 3938
rect 1607 3904 1619 3938
rect 219 3898 352 3904
rect 132 3856 138 3890
rect 172 3856 178 3890
rect 342 3888 352 3898
rect 858 3898 1619 3904
rect 858 3888 868 3898
rect 132 3698 178 3856
rect 970 3848 980 3858
rect 219 3842 980 3848
rect 1490 3848 1500 3858
rect 1490 3842 1619 3848
rect 219 3808 231 3842
rect 1607 3808 1619 3842
rect 219 3802 980 3808
rect 970 3792 980 3802
rect 1490 3802 1619 3808
rect 1490 3792 1500 3802
rect 1660 3794 1706 3952
rect 342 3752 352 3762
rect 219 3746 352 3752
rect 858 3752 868 3762
rect 1660 3760 1666 3794
rect 1700 3760 1706 3794
rect 858 3746 1619 3752
rect 219 3712 231 3746
rect 1607 3712 1619 3746
rect 219 3706 352 3712
rect 132 3664 138 3698
rect 172 3664 178 3698
rect 342 3696 352 3706
rect 858 3706 1619 3712
rect 858 3696 868 3706
rect 132 3506 178 3664
rect 970 3656 980 3666
rect 219 3650 980 3656
rect 1490 3656 1500 3666
rect 1490 3650 1619 3656
rect 219 3616 231 3650
rect 1607 3616 1619 3650
rect 219 3610 980 3616
rect 970 3600 980 3610
rect 1490 3610 1619 3616
rect 1490 3600 1500 3610
rect 1660 3602 1706 3760
rect 342 3560 352 3570
rect 219 3554 352 3560
rect 858 3560 868 3570
rect 1660 3568 1666 3602
rect 1700 3568 1706 3602
rect 858 3554 1619 3560
rect 219 3520 231 3554
rect 1607 3520 1619 3554
rect 219 3514 352 3520
rect 132 3472 138 3506
rect 172 3472 178 3506
rect 342 3504 352 3514
rect 858 3514 1619 3520
rect 858 3504 868 3514
rect 132 3314 178 3472
rect 970 3464 980 3474
rect 219 3458 980 3464
rect 1490 3464 1500 3474
rect 1490 3458 1619 3464
rect 219 3424 231 3458
rect 1607 3424 1619 3458
rect 219 3418 980 3424
rect 970 3408 980 3418
rect 1490 3418 1619 3424
rect 1490 3408 1500 3418
rect 1660 3410 1706 3568
rect 342 3368 352 3378
rect 219 3362 352 3368
rect 858 3368 868 3378
rect 1660 3376 1666 3410
rect 1700 3376 1706 3410
rect 858 3362 1619 3368
rect 219 3328 231 3362
rect 1607 3328 1619 3362
rect 219 3322 352 3328
rect 132 3280 138 3314
rect 172 3280 178 3314
rect 342 3312 352 3322
rect 858 3322 1619 3328
rect 858 3312 868 3322
rect 132 3122 178 3280
rect 970 3272 980 3282
rect 219 3266 980 3272
rect 1490 3272 1500 3282
rect 1490 3266 1619 3272
rect 219 3232 231 3266
rect 1607 3232 1619 3266
rect 219 3226 980 3232
rect 970 3216 980 3226
rect 1490 3226 1619 3232
rect 1490 3216 1500 3226
rect 1660 3218 1706 3376
rect 342 3176 352 3186
rect 219 3170 352 3176
rect 858 3176 868 3186
rect 1660 3184 1666 3218
rect 1700 3184 1706 3218
rect 858 3170 1619 3176
rect 219 3136 231 3170
rect 1607 3136 1619 3170
rect 219 3130 352 3136
rect 132 3088 138 3122
rect 172 3088 178 3122
rect 342 3120 352 3130
rect 858 3130 1619 3136
rect 858 3120 868 3130
rect 132 2930 178 3088
rect 970 3080 980 3090
rect 219 3074 980 3080
rect 1490 3080 1500 3090
rect 1490 3074 1619 3080
rect 219 3040 231 3074
rect 1607 3040 1619 3074
rect 219 3034 980 3040
rect 970 3024 980 3034
rect 1490 3034 1619 3040
rect 1490 3024 1500 3034
rect 1660 3026 1706 3184
rect 342 2984 352 2994
rect 219 2978 352 2984
rect 858 2984 868 2994
rect 1660 2992 1666 3026
rect 1700 2992 1706 3026
rect 858 2978 1619 2984
rect 219 2944 231 2978
rect 1607 2944 1619 2978
rect 219 2938 352 2944
rect 132 2896 138 2930
rect 172 2896 178 2930
rect 342 2928 352 2938
rect 858 2938 1619 2944
rect 858 2928 868 2938
rect 132 2738 178 2896
rect 970 2888 980 2898
rect 219 2882 980 2888
rect 1490 2888 1500 2898
rect 1490 2882 1619 2888
rect 219 2848 231 2882
rect 1607 2848 1619 2882
rect 219 2842 980 2848
rect 970 2832 980 2842
rect 1490 2842 1619 2848
rect 1490 2832 1500 2842
rect 1660 2834 1706 2992
rect 342 2792 352 2802
rect 219 2786 352 2792
rect 858 2792 868 2802
rect 1660 2800 1666 2834
rect 1700 2800 1706 2834
rect 858 2786 1619 2792
rect 219 2752 231 2786
rect 1607 2752 1619 2786
rect 219 2746 352 2752
rect 132 2704 138 2738
rect 172 2704 178 2738
rect 342 2736 352 2746
rect 858 2746 1619 2752
rect 858 2736 868 2746
rect 132 2546 178 2704
rect 970 2696 980 2706
rect 219 2690 980 2696
rect 1490 2696 1500 2706
rect 1490 2690 1619 2696
rect 219 2656 231 2690
rect 1607 2656 1619 2690
rect 219 2650 980 2656
rect 970 2640 980 2650
rect 1490 2650 1619 2656
rect 1490 2640 1500 2650
rect 1660 2642 1706 2800
rect 342 2600 352 2610
rect 219 2594 352 2600
rect 858 2600 868 2610
rect 1660 2608 1666 2642
rect 1700 2608 1706 2642
rect 858 2594 1619 2600
rect 219 2560 231 2594
rect 1607 2560 1619 2594
rect 219 2554 352 2560
rect 132 2512 138 2546
rect 172 2512 178 2546
rect 342 2544 352 2554
rect 858 2554 1619 2560
rect 858 2544 868 2554
rect 132 2354 178 2512
rect 970 2504 980 2514
rect 219 2498 980 2504
rect 1490 2504 1500 2514
rect 1490 2498 1619 2504
rect 219 2464 231 2498
rect 1607 2464 1619 2498
rect 219 2458 980 2464
rect 970 2448 980 2458
rect 1490 2458 1619 2464
rect 1490 2448 1500 2458
rect 1660 2450 1706 2608
rect 342 2408 352 2418
rect 219 2402 352 2408
rect 858 2408 868 2418
rect 1660 2416 1666 2450
rect 1700 2416 1706 2450
rect 858 2402 1619 2408
rect 219 2368 231 2402
rect 1607 2368 1619 2402
rect 219 2362 352 2368
rect 132 2320 138 2354
rect 172 2320 178 2354
rect 342 2352 352 2362
rect 858 2362 1619 2368
rect 858 2352 868 2362
rect 132 2162 178 2320
rect 970 2312 980 2322
rect 219 2306 980 2312
rect 1490 2312 1500 2322
rect 1490 2306 1619 2312
rect 219 2272 231 2306
rect 1607 2272 1619 2306
rect 219 2266 980 2272
rect 970 2256 980 2266
rect 1490 2266 1619 2272
rect 1490 2256 1500 2266
rect 1660 2258 1706 2416
rect 342 2216 352 2226
rect 219 2210 352 2216
rect 858 2216 868 2226
rect 1660 2224 1666 2258
rect 1700 2224 1706 2258
rect 858 2210 1619 2216
rect 219 2176 231 2210
rect 1607 2176 1619 2210
rect 219 2170 352 2176
rect 132 2128 138 2162
rect 172 2128 178 2162
rect 342 2160 352 2170
rect 858 2170 1619 2176
rect 858 2160 868 2170
rect 132 1970 178 2128
rect 970 2120 980 2130
rect 219 2114 980 2120
rect 1490 2120 1500 2130
rect 1490 2114 1619 2120
rect 219 2080 231 2114
rect 1607 2080 1619 2114
rect 219 2074 980 2080
rect 970 2064 980 2074
rect 1490 2074 1619 2080
rect 1490 2064 1500 2074
rect 1660 2066 1706 2224
rect 342 2024 352 2034
rect 219 2018 352 2024
rect 858 2024 868 2034
rect 1660 2032 1666 2066
rect 1700 2032 1706 2066
rect 858 2018 1619 2024
rect 219 1984 231 2018
rect 1607 1984 1619 2018
rect 219 1978 352 1984
rect 132 1936 138 1970
rect 172 1936 178 1970
rect 342 1968 352 1978
rect 858 1978 1619 1984
rect 858 1968 868 1978
rect 132 1778 178 1936
rect 970 1928 980 1938
rect 219 1922 980 1928
rect 1490 1928 1500 1938
rect 1490 1922 1619 1928
rect 219 1888 231 1922
rect 1607 1888 1619 1922
rect 219 1882 980 1888
rect 970 1872 980 1882
rect 1490 1882 1619 1888
rect 1490 1872 1500 1882
rect 1660 1874 1706 2032
rect 342 1832 352 1842
rect 219 1826 352 1832
rect 858 1832 868 1842
rect 1660 1840 1666 1874
rect 1700 1840 1706 1874
rect 858 1826 1619 1832
rect 219 1792 231 1826
rect 1607 1792 1619 1826
rect 219 1786 352 1792
rect 132 1744 138 1778
rect 172 1744 178 1778
rect 342 1776 352 1786
rect 858 1786 1619 1792
rect 858 1776 868 1786
rect 132 1586 178 1744
rect 970 1736 980 1746
rect 219 1730 980 1736
rect 1490 1736 1500 1746
rect 1490 1730 1619 1736
rect 219 1696 231 1730
rect 1607 1696 1619 1730
rect 219 1690 980 1696
rect 970 1680 980 1690
rect 1490 1690 1619 1696
rect 1490 1680 1500 1690
rect 1660 1682 1706 1840
rect 342 1640 352 1650
rect 219 1634 352 1640
rect 858 1640 868 1650
rect 1660 1648 1666 1682
rect 1700 1648 1706 1682
rect 858 1634 1619 1640
rect 219 1600 231 1634
rect 1607 1600 1619 1634
rect 219 1594 352 1600
rect 132 1552 138 1586
rect 172 1552 178 1586
rect 342 1584 352 1594
rect 858 1594 1619 1600
rect 858 1584 868 1594
rect 132 1394 178 1552
rect 970 1544 980 1554
rect 219 1538 980 1544
rect 1490 1544 1500 1554
rect 1490 1538 1619 1544
rect 219 1504 231 1538
rect 1607 1504 1619 1538
rect 219 1498 980 1504
rect 970 1488 980 1498
rect 1490 1498 1619 1504
rect 1490 1488 1500 1498
rect 1660 1490 1706 1648
rect 342 1448 352 1458
rect 219 1442 352 1448
rect 858 1448 868 1458
rect 1660 1456 1666 1490
rect 1700 1456 1706 1490
rect 858 1442 1619 1448
rect 219 1408 231 1442
rect 1607 1408 1619 1442
rect 219 1402 352 1408
rect 132 1360 138 1394
rect 172 1360 178 1394
rect 342 1392 352 1402
rect 858 1402 1619 1408
rect 858 1392 868 1402
rect 132 1202 178 1360
rect 970 1352 980 1362
rect 219 1346 980 1352
rect 1490 1352 1500 1362
rect 1490 1346 1619 1352
rect 219 1312 231 1346
rect 1607 1312 1619 1346
rect 219 1306 980 1312
rect 970 1296 980 1306
rect 1490 1306 1619 1312
rect 1490 1296 1500 1306
rect 1660 1298 1706 1456
rect 342 1256 352 1266
rect 219 1250 352 1256
rect 858 1256 868 1266
rect 1660 1264 1666 1298
rect 1700 1264 1706 1298
rect 858 1250 1619 1256
rect 219 1216 231 1250
rect 1607 1216 1619 1250
rect 219 1210 352 1216
rect 132 1168 138 1202
rect 172 1168 178 1202
rect 342 1200 352 1210
rect 858 1210 1619 1216
rect 858 1200 868 1210
rect 132 1010 178 1168
rect 970 1160 980 1170
rect 219 1154 980 1160
rect 1490 1160 1500 1170
rect 1490 1154 1619 1160
rect 219 1120 231 1154
rect 1607 1120 1619 1154
rect 219 1114 980 1120
rect 970 1104 980 1114
rect 1490 1114 1619 1120
rect 1490 1104 1500 1114
rect 1660 1106 1706 1264
rect 342 1064 352 1074
rect 219 1058 352 1064
rect 858 1064 868 1074
rect 1660 1072 1666 1106
rect 1700 1072 1706 1106
rect 858 1058 1619 1064
rect 219 1024 231 1058
rect 1607 1024 1619 1058
rect 219 1018 352 1024
rect 132 976 138 1010
rect 172 976 178 1010
rect 342 1008 352 1018
rect 858 1018 1619 1024
rect 858 1008 868 1018
rect 132 818 178 976
rect 970 968 980 978
rect 219 962 980 968
rect 1490 968 1500 978
rect 1490 962 1619 968
rect 219 928 231 962
rect 1607 928 1619 962
rect 219 922 980 928
rect 970 912 980 922
rect 1490 922 1619 928
rect 1490 912 1500 922
rect 1660 914 1706 1072
rect 342 872 352 882
rect 219 866 352 872
rect 858 872 868 882
rect 1660 880 1666 914
rect 1700 880 1706 914
rect 858 866 1619 872
rect 219 832 231 866
rect 1607 832 1619 866
rect 219 826 352 832
rect 132 784 138 818
rect 172 784 178 818
rect 342 816 352 826
rect 858 826 1619 832
rect 858 816 868 826
rect 132 772 178 784
rect 970 776 980 786
rect 219 770 980 776
rect 1490 776 1500 786
rect 1490 770 1619 776
rect 219 736 231 770
rect 1607 736 1619 770
rect 219 730 980 736
rect 970 720 980 730
rect 1490 730 1619 736
rect 1490 720 1500 730
rect 1660 722 1706 880
rect 342 680 352 690
rect 219 674 352 680
rect 858 680 868 690
rect 1660 688 1666 722
rect 1700 688 1706 722
rect 858 674 1619 680
rect 1660 676 1706 688
rect 219 640 231 674
rect 1607 640 1619 674
rect 219 634 352 640
rect 342 624 352 634
rect 858 634 1619 640
rect 858 624 868 634
<< via1 >>
rect 132 22222 1706 22286
rect 352 21932 858 21934
rect 342 21868 868 21932
rect 352 21794 858 21810
rect 352 21760 858 21794
rect 352 21744 858 21760
rect 980 21698 1490 21714
rect 980 21664 1490 21698
rect 980 21648 1490 21664
rect 352 21602 858 21618
rect 352 21568 858 21602
rect 352 21552 858 21568
rect 980 21506 1490 21522
rect 980 21472 1490 21506
rect 980 21456 1490 21472
rect 352 21410 858 21426
rect 352 21376 858 21410
rect 352 21360 858 21376
rect 980 21314 1490 21330
rect 980 21280 1490 21314
rect 980 21264 1490 21280
rect 352 21218 858 21234
rect 352 21184 858 21218
rect 352 21168 858 21184
rect 980 21122 1490 21138
rect 980 21088 1490 21122
rect 980 21072 1490 21088
rect 352 21026 858 21042
rect 352 20992 858 21026
rect 352 20976 858 20992
rect 980 20930 1490 20946
rect 980 20896 1490 20930
rect 980 20880 1490 20896
rect 352 20834 858 20850
rect 352 20800 858 20834
rect 352 20784 858 20800
rect 980 20738 1490 20754
rect 980 20704 1490 20738
rect 980 20688 1490 20704
rect 352 20642 858 20658
rect 352 20608 858 20642
rect 352 20592 858 20608
rect 980 20546 1490 20562
rect 980 20512 1490 20546
rect 980 20496 1490 20512
rect 352 20450 858 20466
rect 352 20416 858 20450
rect 352 20400 858 20416
rect 980 20354 1490 20370
rect 980 20320 1490 20354
rect 980 20304 1490 20320
rect 352 20258 858 20274
rect 352 20224 858 20258
rect 352 20208 858 20224
rect 980 20162 1490 20178
rect 980 20128 1490 20162
rect 980 20112 1490 20128
rect 352 20066 858 20082
rect 352 20032 858 20066
rect 352 20016 858 20032
rect 980 19970 1490 19986
rect 980 19936 1490 19970
rect 980 19920 1490 19936
rect 352 19874 858 19890
rect 352 19840 858 19874
rect 352 19824 858 19840
rect 980 19778 1490 19794
rect 980 19744 1490 19778
rect 980 19728 1490 19744
rect 352 19682 858 19698
rect 352 19648 858 19682
rect 352 19632 858 19648
rect 980 19586 1490 19602
rect 980 19552 1490 19586
rect 980 19536 1490 19552
rect 352 19490 858 19506
rect 352 19456 858 19490
rect 352 19440 858 19456
rect 980 19394 1490 19410
rect 980 19360 1490 19394
rect 980 19344 1490 19360
rect 352 19298 858 19314
rect 352 19264 858 19298
rect 352 19248 858 19264
rect 980 19202 1490 19218
rect 980 19168 1490 19202
rect 980 19152 1490 19168
rect 352 19106 858 19122
rect 352 19072 858 19106
rect 352 19056 858 19072
rect 980 19010 1490 19026
rect 980 18976 1490 19010
rect 980 18960 1490 18976
rect 352 18914 858 18930
rect 352 18880 858 18914
rect 352 18864 858 18880
rect 980 18818 1490 18834
rect 980 18784 1490 18818
rect 980 18768 1490 18784
rect 352 18722 858 18738
rect 352 18688 858 18722
rect 352 18672 858 18688
rect 980 18626 1490 18642
rect 980 18592 1490 18626
rect 980 18576 1490 18592
rect 352 18530 858 18546
rect 352 18496 858 18530
rect 352 18480 858 18496
rect 980 18434 1490 18450
rect 980 18400 1490 18434
rect 980 18384 1490 18400
rect 352 18338 858 18354
rect 352 18304 858 18338
rect 352 18288 858 18304
rect 980 18242 1490 18258
rect 980 18208 1490 18242
rect 980 18192 1490 18208
rect 352 18146 858 18162
rect 352 18112 858 18146
rect 352 18096 858 18112
rect 980 18050 1490 18066
rect 980 18016 1490 18050
rect 980 18000 1490 18016
rect 352 17954 858 17970
rect 352 17920 858 17954
rect 352 17904 858 17920
rect 980 17858 1490 17874
rect 980 17824 1490 17858
rect 980 17808 1490 17824
rect 352 17762 858 17778
rect 352 17728 858 17762
rect 352 17712 858 17728
rect 980 17666 1490 17682
rect 980 17632 1490 17666
rect 980 17616 1490 17632
rect 352 17570 858 17586
rect 352 17536 858 17570
rect 352 17520 858 17536
rect 980 17474 1490 17490
rect 980 17440 1490 17474
rect 980 17424 1490 17440
rect 352 17378 858 17394
rect 352 17344 858 17378
rect 352 17328 858 17344
rect 980 17282 1490 17298
rect 980 17248 1490 17282
rect 980 17232 1490 17248
rect 352 17186 858 17202
rect 352 17152 858 17186
rect 352 17136 858 17152
rect 980 17090 1490 17106
rect 980 17056 1490 17090
rect 980 17040 1490 17056
rect 352 16994 858 17010
rect 352 16960 858 16994
rect 352 16944 858 16960
rect 980 16898 1490 16914
rect 980 16864 1490 16898
rect 980 16848 1490 16864
rect 352 16802 858 16818
rect 352 16768 858 16802
rect 352 16752 858 16768
rect 980 16706 1490 16722
rect 980 16672 1490 16706
rect 980 16656 1490 16672
rect 352 16610 858 16626
rect 352 16576 858 16610
rect 352 16560 858 16576
rect 980 16514 1490 16530
rect 980 16480 1490 16514
rect 980 16464 1490 16480
rect 352 16418 858 16434
rect 352 16384 858 16418
rect 352 16368 858 16384
rect 980 16322 1490 16338
rect 980 16288 1490 16322
rect 980 16272 1490 16288
rect 352 16226 858 16242
rect 352 16192 858 16226
rect 352 16176 858 16192
rect 980 16130 1490 16146
rect 980 16096 1490 16130
rect 980 16080 1490 16096
rect 352 16034 858 16050
rect 352 16000 858 16034
rect 352 15984 858 16000
rect 980 15938 1490 15954
rect 980 15904 1490 15938
rect 980 15888 1490 15904
rect 352 15842 858 15858
rect 352 15808 858 15842
rect 352 15792 858 15808
rect 980 15746 1490 15762
rect 980 15712 1490 15746
rect 980 15696 1490 15712
rect 352 15650 858 15666
rect 352 15616 858 15650
rect 352 15600 858 15616
rect 980 15554 1490 15570
rect 980 15520 1490 15554
rect 980 15504 1490 15520
rect 352 15458 858 15474
rect 352 15424 858 15458
rect 352 15408 858 15424
rect 980 15362 1490 15378
rect 980 15328 1490 15362
rect 980 15312 1490 15328
rect 352 15266 858 15282
rect 352 15232 858 15266
rect 352 15216 858 15232
rect 980 15170 1490 15186
rect 980 15136 1490 15170
rect 980 15120 1490 15136
rect 352 15074 858 15090
rect 352 15040 858 15074
rect 352 15024 858 15040
rect 980 14978 1490 14994
rect 980 14944 1490 14978
rect 980 14928 1490 14944
rect 352 14882 858 14898
rect 352 14848 858 14882
rect 352 14832 858 14848
rect 980 14786 1490 14802
rect 980 14752 1490 14786
rect 980 14736 1490 14752
rect 352 14690 858 14706
rect 352 14656 858 14690
rect 352 14640 858 14656
rect 980 14594 1490 14610
rect 980 14560 1490 14594
rect 980 14544 1490 14560
rect 352 14498 858 14514
rect 352 14464 858 14498
rect 352 14448 858 14464
rect 980 14402 1490 14418
rect 980 14368 1490 14402
rect 980 14352 1490 14368
rect 352 14306 858 14322
rect 352 14272 858 14306
rect 352 14256 858 14272
rect 980 14210 1490 14226
rect 980 14176 1490 14210
rect 980 14160 1490 14176
rect 352 14114 858 14130
rect 352 14080 858 14114
rect 352 14064 858 14080
rect 980 14018 1490 14034
rect 980 13984 1490 14018
rect 980 13968 1490 13984
rect 352 13922 858 13938
rect 352 13888 858 13922
rect 352 13872 858 13888
rect 980 13826 1490 13842
rect 980 13792 1490 13826
rect 980 13776 1490 13792
rect 352 13730 858 13746
rect 352 13696 858 13730
rect 352 13680 858 13696
rect 980 13634 1490 13650
rect 980 13600 1490 13634
rect 980 13584 1490 13600
rect 352 13538 858 13554
rect 352 13504 858 13538
rect 352 13488 858 13504
rect 980 13442 1490 13458
rect 980 13408 1490 13442
rect 980 13392 1490 13408
rect 352 13346 858 13362
rect 352 13312 858 13346
rect 352 13296 858 13312
rect 980 13250 1490 13266
rect 980 13216 1490 13250
rect 980 13200 1490 13216
rect 352 13154 858 13170
rect 352 13120 858 13154
rect 352 13104 858 13120
rect 980 13058 1490 13074
rect 980 13024 1490 13058
rect 980 13008 1490 13024
rect 352 12962 858 12978
rect 352 12928 858 12962
rect 352 12912 858 12928
rect 980 12866 1490 12882
rect 980 12832 1490 12866
rect 980 12816 1490 12832
rect 352 12770 858 12786
rect 352 12736 858 12770
rect 352 12720 858 12736
rect 980 12674 1490 12690
rect 980 12640 1490 12674
rect 980 12624 1490 12640
rect 352 12578 858 12594
rect 352 12544 858 12578
rect 352 12528 858 12544
rect 980 12482 1490 12498
rect 980 12448 1490 12482
rect 980 12432 1490 12448
rect 352 12386 858 12402
rect 352 12352 858 12386
rect 352 12336 858 12352
rect 980 12290 1490 12306
rect 980 12256 1490 12290
rect 980 12240 1490 12256
rect 352 12194 858 12210
rect 352 12160 858 12194
rect 352 12144 858 12160
rect 980 12098 1490 12114
rect 980 12064 1490 12098
rect 980 12048 1490 12064
rect 352 12002 858 12018
rect 352 11968 858 12002
rect 352 11952 858 11968
rect 980 11906 1490 11922
rect 980 11872 1490 11906
rect 980 11856 1490 11872
rect 352 11810 858 11826
rect 352 11776 858 11810
rect 352 11760 858 11776
rect 980 11714 1490 11730
rect 980 11680 1490 11714
rect 980 11664 1490 11680
rect 352 11618 858 11634
rect 352 11584 858 11618
rect 352 11568 858 11584
rect 980 11522 1490 11538
rect 980 11488 1490 11522
rect 980 11472 1490 11488
rect 352 11426 858 11442
rect 352 11392 858 11426
rect 352 11376 858 11392
rect 980 11330 1490 11346
rect 980 11296 1490 11330
rect 980 11280 1490 11296
rect 352 11234 858 11250
rect 352 11200 858 11234
rect 352 11184 858 11200
rect 980 11138 1490 11154
rect 980 11104 1490 11138
rect 980 11088 1490 11104
rect 352 11042 858 11058
rect 352 11008 858 11042
rect 352 10992 858 11008
rect 980 10946 1490 10962
rect 980 10912 1490 10946
rect 980 10896 1490 10912
rect 352 10850 858 10866
rect 352 10816 858 10850
rect 352 10800 858 10816
rect 980 10754 1490 10770
rect 980 10720 1490 10754
rect 980 10704 1490 10720
rect 352 10658 858 10674
rect 352 10624 858 10658
rect 352 10608 858 10624
rect 980 10562 1490 10578
rect 980 10528 1490 10562
rect 980 10512 1490 10528
rect 352 10466 858 10482
rect 352 10432 858 10466
rect 352 10416 858 10432
rect 980 10370 1490 10386
rect 980 10336 1490 10370
rect 980 10320 1490 10336
rect 352 10274 858 10290
rect 352 10240 858 10274
rect 352 10224 858 10240
rect 980 10178 1490 10194
rect 980 10144 1490 10178
rect 980 10128 1490 10144
rect 352 10082 858 10098
rect 352 10048 858 10082
rect 352 10032 858 10048
rect 980 9986 1490 10002
rect 980 9952 1490 9986
rect 980 9936 1490 9952
rect 352 9890 858 9906
rect 352 9856 858 9890
rect 352 9840 858 9856
rect 980 9794 1490 9810
rect 980 9760 1490 9794
rect 980 9744 1490 9760
rect 352 9698 858 9714
rect 352 9664 858 9698
rect 352 9648 858 9664
rect 980 9602 1490 9618
rect 980 9568 1490 9602
rect 980 9552 1490 9568
rect 352 9506 858 9522
rect 352 9472 858 9506
rect 352 9456 858 9472
rect 980 9410 1490 9426
rect 980 9376 1490 9410
rect 980 9360 1490 9376
rect 352 9314 858 9330
rect 352 9280 858 9314
rect 352 9264 858 9280
rect 980 9218 1490 9234
rect 980 9184 1490 9218
rect 980 9168 1490 9184
rect 352 9122 858 9138
rect 352 9088 858 9122
rect 352 9072 858 9088
rect 980 9026 1490 9042
rect 980 8992 1490 9026
rect 980 8976 1490 8992
rect 352 8930 858 8946
rect 352 8896 858 8930
rect 352 8880 858 8896
rect 980 8834 1490 8850
rect 980 8800 1490 8834
rect 980 8784 1490 8800
rect 352 8738 858 8754
rect 352 8704 858 8738
rect 352 8688 858 8704
rect 980 8642 1490 8658
rect 980 8608 1490 8642
rect 980 8592 1490 8608
rect 352 8546 858 8562
rect 352 8512 858 8546
rect 352 8496 858 8512
rect 980 8450 1490 8466
rect 980 8416 1490 8450
rect 980 8400 1490 8416
rect 352 8354 858 8370
rect 352 8320 858 8354
rect 352 8304 858 8320
rect 980 8258 1490 8274
rect 980 8224 1490 8258
rect 980 8208 1490 8224
rect 352 8162 858 8178
rect 352 8128 858 8162
rect 352 8112 858 8128
rect 980 8066 1490 8082
rect 980 8032 1490 8066
rect 980 8016 1490 8032
rect 352 7970 858 7986
rect 352 7936 858 7970
rect 352 7920 858 7936
rect 980 7874 1490 7890
rect 980 7840 1490 7874
rect 980 7824 1490 7840
rect 352 7778 858 7794
rect 352 7744 858 7778
rect 352 7728 858 7744
rect 980 7682 1490 7698
rect 980 7648 1490 7682
rect 980 7632 1490 7648
rect 352 7586 858 7602
rect 352 7552 858 7586
rect 352 7536 858 7552
rect 980 7490 1490 7506
rect 980 7456 1490 7490
rect 980 7440 1490 7456
rect 352 7394 858 7410
rect 352 7360 858 7394
rect 352 7344 858 7360
rect 980 7298 1490 7314
rect 980 7264 1490 7298
rect 980 7248 1490 7264
rect 352 7202 858 7218
rect 352 7168 858 7202
rect 352 7152 858 7168
rect 980 7106 1490 7122
rect 980 7072 1490 7106
rect 980 7056 1490 7072
rect 352 7010 858 7026
rect 352 6976 858 7010
rect 352 6960 858 6976
rect 980 6914 1490 6930
rect 980 6880 1490 6914
rect 980 6864 1490 6880
rect 352 6818 858 6834
rect 352 6784 858 6818
rect 352 6768 858 6784
rect 980 6722 1490 6738
rect 980 6688 1490 6722
rect 980 6672 1490 6688
rect 352 6626 858 6642
rect 352 6592 858 6626
rect 352 6576 858 6592
rect 980 6530 1490 6546
rect 980 6496 1490 6530
rect 980 6480 1490 6496
rect 352 6434 858 6450
rect 352 6400 858 6434
rect 352 6384 858 6400
rect 980 6338 1490 6354
rect 980 6304 1490 6338
rect 980 6288 1490 6304
rect 352 6242 858 6258
rect 352 6208 858 6242
rect 352 6192 858 6208
rect 980 6146 1490 6162
rect 980 6112 1490 6146
rect 980 6096 1490 6112
rect 352 6050 858 6066
rect 352 6016 858 6050
rect 352 6000 858 6016
rect 980 5954 1490 5970
rect 980 5920 1490 5954
rect 980 5904 1490 5920
rect 352 5858 858 5874
rect 352 5824 858 5858
rect 352 5808 858 5824
rect 980 5762 1490 5778
rect 980 5728 1490 5762
rect 980 5712 1490 5728
rect 352 5666 858 5682
rect 352 5632 858 5666
rect 352 5616 858 5632
rect 980 5570 1490 5586
rect 980 5536 1490 5570
rect 980 5520 1490 5536
rect 352 5474 858 5490
rect 352 5440 858 5474
rect 352 5424 858 5440
rect 980 5378 1490 5394
rect 980 5344 1490 5378
rect 980 5328 1490 5344
rect 352 5282 858 5298
rect 352 5248 858 5282
rect 352 5232 858 5248
rect 980 5186 1490 5202
rect 980 5152 1490 5186
rect 980 5136 1490 5152
rect 352 5090 858 5106
rect 352 5056 858 5090
rect 352 5040 858 5056
rect 980 4994 1490 5010
rect 980 4960 1490 4994
rect 980 4944 1490 4960
rect 352 4898 858 4914
rect 352 4864 858 4898
rect 352 4848 858 4864
rect 980 4802 1490 4818
rect 980 4768 1490 4802
rect 980 4752 1490 4768
rect 352 4706 858 4722
rect 352 4672 858 4706
rect 352 4656 858 4672
rect 980 4610 1490 4626
rect 980 4576 1490 4610
rect 980 4560 1490 4576
rect 352 4514 858 4530
rect 352 4480 858 4514
rect 352 4464 858 4480
rect 980 4418 1490 4434
rect 980 4384 1490 4418
rect 980 4368 1490 4384
rect 352 4322 858 4338
rect 352 4288 858 4322
rect 352 4272 858 4288
rect 980 4226 1490 4242
rect 980 4192 1490 4226
rect 980 4176 1490 4192
rect 352 4130 858 4146
rect 352 4096 858 4130
rect 352 4080 858 4096
rect 980 4034 1490 4050
rect 980 4000 1490 4034
rect 980 3984 1490 4000
rect 352 3938 858 3954
rect 352 3904 858 3938
rect 352 3888 858 3904
rect 980 3842 1490 3858
rect 980 3808 1490 3842
rect 980 3792 1490 3808
rect 352 3746 858 3762
rect 352 3712 858 3746
rect 352 3696 858 3712
rect 980 3650 1490 3666
rect 980 3616 1490 3650
rect 980 3600 1490 3616
rect 352 3554 858 3570
rect 352 3520 858 3554
rect 352 3504 858 3520
rect 980 3458 1490 3474
rect 980 3424 1490 3458
rect 980 3408 1490 3424
rect 352 3362 858 3378
rect 352 3328 858 3362
rect 352 3312 858 3328
rect 980 3266 1490 3282
rect 980 3232 1490 3266
rect 980 3216 1490 3232
rect 352 3170 858 3186
rect 352 3136 858 3170
rect 352 3120 858 3136
rect 980 3074 1490 3090
rect 980 3040 1490 3074
rect 980 3024 1490 3040
rect 352 2978 858 2994
rect 352 2944 858 2978
rect 352 2928 858 2944
rect 980 2882 1490 2898
rect 980 2848 1490 2882
rect 980 2832 1490 2848
rect 352 2786 858 2802
rect 352 2752 858 2786
rect 352 2736 858 2752
rect 980 2690 1490 2706
rect 980 2656 1490 2690
rect 980 2640 1490 2656
rect 352 2594 858 2610
rect 352 2560 858 2594
rect 352 2544 858 2560
rect 980 2498 1490 2514
rect 980 2464 1490 2498
rect 980 2448 1490 2464
rect 352 2402 858 2418
rect 352 2368 858 2402
rect 352 2352 858 2368
rect 980 2306 1490 2322
rect 980 2272 1490 2306
rect 980 2256 1490 2272
rect 352 2210 858 2226
rect 352 2176 858 2210
rect 352 2160 858 2176
rect 980 2114 1490 2130
rect 980 2080 1490 2114
rect 980 2064 1490 2080
rect 352 2018 858 2034
rect 352 1984 858 2018
rect 352 1968 858 1984
rect 980 1922 1490 1938
rect 980 1888 1490 1922
rect 980 1872 1490 1888
rect 352 1826 858 1842
rect 352 1792 858 1826
rect 352 1776 858 1792
rect 980 1730 1490 1746
rect 980 1696 1490 1730
rect 980 1680 1490 1696
rect 352 1634 858 1650
rect 352 1600 858 1634
rect 352 1584 858 1600
rect 980 1538 1490 1554
rect 980 1504 1490 1538
rect 980 1488 1490 1504
rect 352 1442 858 1458
rect 352 1408 858 1442
rect 352 1392 858 1408
rect 980 1346 1490 1362
rect 980 1312 1490 1346
rect 980 1296 1490 1312
rect 352 1250 858 1266
rect 352 1216 858 1250
rect 352 1200 858 1216
rect 980 1154 1490 1170
rect 980 1120 1490 1154
rect 980 1104 1490 1120
rect 352 1058 858 1074
rect 352 1024 858 1058
rect 352 1008 858 1024
rect 980 962 1490 978
rect 980 928 1490 962
rect 980 912 1490 928
rect 352 866 858 882
rect 352 832 858 866
rect 352 816 858 832
rect 980 770 1490 786
rect 980 736 1490 770
rect 980 720 1490 736
rect 352 674 858 690
rect 352 640 858 674
rect 352 624 858 640
<< metal2 >>
rect 132 22286 1706 22296
rect 132 22212 1706 22222
rect 342 21934 868 21942
rect 342 21932 352 21934
rect 858 21932 868 21934
rect 342 21858 868 21868
rect 342 21810 868 21820
rect 342 21744 352 21810
rect 858 21744 868 21810
rect 342 21734 868 21744
rect 970 21714 1500 21724
rect 970 21648 980 21714
rect 1490 21648 1500 21714
rect 970 21638 1500 21648
rect 342 21618 868 21628
rect 342 21552 352 21618
rect 858 21552 868 21618
rect 342 21542 868 21552
rect 970 21522 1500 21532
rect 970 21456 980 21522
rect 1490 21456 1500 21522
rect 970 21446 1500 21456
rect 342 21426 868 21436
rect 342 21360 352 21426
rect 858 21360 868 21426
rect 342 21350 868 21360
rect 970 21330 1500 21340
rect 970 21264 980 21330
rect 1490 21264 1500 21330
rect 970 21254 1500 21264
rect 342 21234 868 21244
rect 342 21168 352 21234
rect 858 21168 868 21234
rect 342 21158 868 21168
rect 970 21138 1500 21148
rect 970 21072 980 21138
rect 1490 21072 1500 21138
rect 970 21062 1500 21072
rect 342 21042 868 21052
rect 342 20976 352 21042
rect 858 20976 868 21042
rect 342 20966 868 20976
rect 970 20946 1500 20956
rect 970 20880 980 20946
rect 1490 20880 1500 20946
rect 970 20870 1500 20880
rect 342 20850 868 20860
rect 342 20784 352 20850
rect 858 20784 868 20850
rect 342 20774 868 20784
rect 970 20754 1500 20764
rect 970 20688 980 20754
rect 1490 20688 1500 20754
rect 970 20678 1500 20688
rect 342 20658 868 20668
rect 342 20592 352 20658
rect 858 20592 868 20658
rect 342 20582 868 20592
rect 970 20562 1500 20572
rect 970 20496 980 20562
rect 1490 20496 1500 20562
rect 970 20486 1500 20496
rect 342 20466 868 20476
rect 342 20400 352 20466
rect 858 20400 868 20466
rect 342 20390 868 20400
rect 970 20370 1500 20380
rect 970 20304 980 20370
rect 1490 20304 1500 20370
rect 970 20294 1500 20304
rect 342 20274 868 20284
rect 342 20208 352 20274
rect 858 20208 868 20274
rect 342 20198 868 20208
rect 970 20178 1500 20188
rect 970 20112 980 20178
rect 1490 20112 1500 20178
rect 970 20102 1500 20112
rect 342 20082 868 20092
rect 342 20016 352 20082
rect 858 20016 868 20082
rect 342 20006 868 20016
rect 970 19986 1500 19996
rect 970 19920 980 19986
rect 1490 19920 1500 19986
rect 970 19910 1500 19920
rect 342 19890 868 19900
rect 342 19824 352 19890
rect 858 19824 868 19890
rect 342 19814 868 19824
rect 970 19794 1500 19804
rect 970 19728 980 19794
rect 1490 19728 1500 19794
rect 970 19718 1500 19728
rect 342 19698 868 19708
rect 342 19632 352 19698
rect 858 19632 868 19698
rect 342 19622 868 19632
rect 970 19602 1500 19612
rect 970 19536 980 19602
rect 1490 19536 1500 19602
rect 970 19526 1500 19536
rect 342 19506 868 19516
rect 342 19440 352 19506
rect 858 19440 868 19506
rect 342 19430 868 19440
rect 970 19410 1500 19420
rect 970 19344 980 19410
rect 1490 19344 1500 19410
rect 970 19334 1500 19344
rect 342 19314 868 19324
rect 342 19248 352 19314
rect 858 19248 868 19314
rect 342 19238 868 19248
rect 970 19218 1500 19228
rect 970 19152 980 19218
rect 1490 19152 1500 19218
rect 970 19142 1500 19152
rect 342 19122 868 19132
rect 342 19056 352 19122
rect 858 19056 868 19122
rect 342 19046 868 19056
rect 970 19026 1500 19036
rect 970 18960 980 19026
rect 1490 18960 1500 19026
rect 970 18950 1500 18960
rect 342 18930 868 18940
rect 342 18864 352 18930
rect 858 18864 868 18930
rect 342 18854 868 18864
rect 970 18834 1500 18844
rect 970 18768 980 18834
rect 1490 18768 1500 18834
rect 970 18758 1500 18768
rect 342 18738 868 18748
rect 342 18672 352 18738
rect 858 18672 868 18738
rect 342 18662 868 18672
rect 970 18642 1500 18652
rect 970 18576 980 18642
rect 1490 18576 1500 18642
rect 970 18566 1500 18576
rect 342 18546 868 18556
rect 342 18480 352 18546
rect 858 18480 868 18546
rect 342 18470 868 18480
rect 970 18450 1500 18460
rect 970 18384 980 18450
rect 1490 18384 1500 18450
rect 970 18374 1500 18384
rect 342 18354 868 18364
rect 342 18288 352 18354
rect 858 18288 868 18354
rect 342 18278 868 18288
rect 970 18258 1500 18268
rect 970 18192 980 18258
rect 1490 18192 1500 18258
rect 970 18182 1500 18192
rect 342 18162 868 18172
rect 342 18096 352 18162
rect 858 18096 868 18162
rect 342 18086 868 18096
rect 970 18066 1500 18076
rect 970 18000 980 18066
rect 1490 18000 1500 18066
rect 970 17990 1500 18000
rect 342 17970 868 17980
rect 342 17904 352 17970
rect 858 17904 868 17970
rect 342 17894 868 17904
rect 970 17874 1500 17884
rect 970 17808 980 17874
rect 1490 17808 1500 17874
rect 970 17798 1500 17808
rect 342 17778 868 17788
rect 342 17712 352 17778
rect 858 17712 868 17778
rect 342 17702 868 17712
rect 970 17682 1500 17692
rect 970 17616 980 17682
rect 1490 17616 1500 17682
rect 970 17606 1500 17616
rect 342 17586 868 17596
rect 342 17520 352 17586
rect 858 17520 868 17586
rect 342 17510 868 17520
rect 970 17490 1500 17500
rect 970 17424 980 17490
rect 1490 17424 1500 17490
rect 970 17414 1500 17424
rect 342 17394 868 17404
rect 342 17328 352 17394
rect 858 17328 868 17394
rect 342 17318 868 17328
rect 970 17298 1500 17308
rect 970 17232 980 17298
rect 1490 17232 1500 17298
rect 970 17222 1500 17232
rect 342 17202 868 17212
rect 342 17136 352 17202
rect 858 17136 868 17202
rect 342 17126 868 17136
rect 970 17106 1500 17116
rect 970 17040 980 17106
rect 1490 17040 1500 17106
rect 970 17030 1500 17040
rect 342 17010 868 17020
rect 342 16944 352 17010
rect 858 16944 868 17010
rect 342 16934 868 16944
rect 970 16914 1500 16924
rect 970 16848 980 16914
rect 1490 16848 1500 16914
rect 970 16838 1500 16848
rect 342 16818 868 16828
rect 342 16752 352 16818
rect 858 16752 868 16818
rect 342 16742 868 16752
rect 970 16722 1500 16732
rect 970 16656 980 16722
rect 1490 16656 1500 16722
rect 970 16646 1500 16656
rect 342 16626 868 16636
rect 342 16560 352 16626
rect 858 16560 868 16626
rect 342 16550 868 16560
rect 970 16530 1500 16540
rect 970 16464 980 16530
rect 1490 16464 1500 16530
rect 970 16454 1500 16464
rect 342 16434 868 16444
rect 342 16368 352 16434
rect 858 16368 868 16434
rect 342 16358 868 16368
rect 970 16338 1500 16348
rect 970 16272 980 16338
rect 1490 16272 1500 16338
rect 970 16262 1500 16272
rect 342 16242 868 16252
rect 342 16176 352 16242
rect 858 16176 868 16242
rect 342 16166 868 16176
rect 970 16146 1500 16156
rect 970 16080 980 16146
rect 1490 16080 1500 16146
rect 970 16070 1500 16080
rect 342 16050 868 16060
rect 342 15984 352 16050
rect 858 15984 868 16050
rect 342 15974 868 15984
rect 970 15954 1500 15964
rect 970 15888 980 15954
rect 1490 15888 1500 15954
rect 970 15878 1500 15888
rect 342 15858 868 15868
rect 342 15792 352 15858
rect 858 15792 868 15858
rect 342 15782 868 15792
rect 970 15762 1500 15772
rect 970 15696 980 15762
rect 1490 15696 1500 15762
rect 970 15686 1500 15696
rect 342 15666 868 15676
rect 342 15600 352 15666
rect 858 15600 868 15666
rect 342 15590 868 15600
rect 970 15570 1500 15580
rect 970 15504 980 15570
rect 1490 15504 1500 15570
rect 970 15494 1500 15504
rect 342 15474 868 15484
rect 342 15408 352 15474
rect 858 15408 868 15474
rect 342 15398 868 15408
rect 970 15378 1500 15388
rect 970 15312 980 15378
rect 1490 15312 1500 15378
rect 970 15302 1500 15312
rect 342 15282 868 15292
rect 342 15216 352 15282
rect 858 15216 868 15282
rect 342 15206 868 15216
rect 970 15186 1500 15196
rect 970 15120 980 15186
rect 1490 15120 1500 15186
rect 970 15110 1500 15120
rect 342 15090 868 15100
rect 342 15024 352 15090
rect 858 15024 868 15090
rect 342 15014 868 15024
rect 970 14994 1500 15004
rect 970 14928 980 14994
rect 1490 14928 1500 14994
rect 970 14918 1500 14928
rect 342 14898 868 14908
rect 342 14832 352 14898
rect 858 14832 868 14898
rect 342 14822 868 14832
rect 970 14802 1500 14812
rect 970 14736 980 14802
rect 1490 14736 1500 14802
rect 970 14726 1500 14736
rect 342 14706 868 14716
rect 342 14640 352 14706
rect 858 14640 868 14706
rect 342 14630 868 14640
rect 970 14610 1500 14620
rect 970 14544 980 14610
rect 1490 14544 1500 14610
rect 970 14534 1500 14544
rect 342 14514 868 14524
rect 342 14448 352 14514
rect 858 14448 868 14514
rect 342 14438 868 14448
rect 970 14418 1500 14428
rect 970 14352 980 14418
rect 1490 14352 1500 14418
rect 970 14342 1500 14352
rect 342 14322 868 14332
rect 342 14256 352 14322
rect 858 14256 868 14322
rect 342 14246 868 14256
rect 970 14226 1500 14236
rect 970 14160 980 14226
rect 1490 14160 1500 14226
rect 970 14150 1500 14160
rect 342 14130 868 14140
rect 342 14064 352 14130
rect 858 14064 868 14130
rect 342 14054 868 14064
rect 970 14034 1500 14044
rect 970 13968 980 14034
rect 1490 13968 1500 14034
rect 970 13958 1500 13968
rect 342 13938 868 13948
rect 342 13872 352 13938
rect 858 13872 868 13938
rect 342 13862 868 13872
rect 970 13842 1500 13852
rect 970 13776 980 13842
rect 1490 13776 1500 13842
rect 970 13766 1500 13776
rect 342 13746 868 13756
rect 342 13680 352 13746
rect 858 13680 868 13746
rect 342 13670 868 13680
rect 970 13650 1500 13660
rect 970 13584 980 13650
rect 1490 13584 1500 13650
rect 970 13574 1500 13584
rect 342 13554 868 13564
rect 342 13488 352 13554
rect 858 13488 868 13554
rect 342 13478 868 13488
rect 970 13458 1500 13468
rect 970 13392 980 13458
rect 1490 13392 1500 13458
rect 970 13382 1500 13392
rect 342 13362 868 13372
rect 342 13296 352 13362
rect 858 13296 868 13362
rect 342 13286 868 13296
rect 970 13266 1500 13276
rect 970 13200 980 13266
rect 1490 13200 1500 13266
rect 970 13190 1500 13200
rect 342 13170 868 13180
rect 342 13104 352 13170
rect 858 13104 868 13170
rect 342 13094 868 13104
rect 970 13074 1500 13084
rect 970 13008 980 13074
rect 1490 13008 1500 13074
rect 970 12998 1500 13008
rect 342 12978 868 12988
rect 342 12912 352 12978
rect 858 12912 868 12978
rect 342 12902 868 12912
rect 970 12882 1500 12892
rect 970 12816 980 12882
rect 1490 12816 1500 12882
rect 970 12806 1500 12816
rect 342 12786 868 12796
rect 342 12720 352 12786
rect 858 12720 868 12786
rect 342 12710 868 12720
rect 970 12690 1500 12700
rect 970 12624 980 12690
rect 1490 12624 1500 12690
rect 970 12614 1500 12624
rect 342 12594 868 12604
rect 342 12528 352 12594
rect 858 12528 868 12594
rect 342 12518 868 12528
rect 970 12498 1500 12508
rect 970 12432 980 12498
rect 1490 12432 1500 12498
rect 970 12422 1500 12432
rect 342 12402 868 12412
rect 342 12336 352 12402
rect 858 12336 868 12402
rect 342 12326 868 12336
rect 970 12306 1500 12316
rect 970 12240 980 12306
rect 1490 12240 1500 12306
rect 970 12230 1500 12240
rect 342 12210 868 12220
rect 342 12144 352 12210
rect 858 12144 868 12210
rect 342 12134 868 12144
rect 970 12114 1500 12124
rect 970 12048 980 12114
rect 1490 12048 1500 12114
rect 970 12038 1500 12048
rect 342 12018 868 12028
rect 342 11952 352 12018
rect 858 11952 868 12018
rect 342 11942 868 11952
rect 970 11922 1500 11932
rect 970 11856 980 11922
rect 1490 11856 1500 11922
rect 970 11846 1500 11856
rect 342 11826 868 11836
rect 342 11760 352 11826
rect 858 11760 868 11826
rect 342 11750 868 11760
rect 970 11730 1500 11740
rect 970 11664 980 11730
rect 1490 11664 1500 11730
rect 970 11654 1500 11664
rect 342 11634 868 11644
rect 342 11568 352 11634
rect 858 11568 868 11634
rect 342 11558 868 11568
rect 970 11538 1500 11548
rect 970 11472 980 11538
rect 1490 11472 1500 11538
rect 970 11462 1500 11472
rect 342 11442 868 11452
rect 342 11376 352 11442
rect 858 11376 868 11442
rect 342 11366 868 11376
rect 970 11346 1500 11356
rect 970 11280 980 11346
rect 1490 11280 1500 11346
rect 970 11270 1500 11280
rect 342 11250 868 11260
rect 342 11184 352 11250
rect 858 11184 868 11250
rect 342 11174 868 11184
rect 970 11154 1500 11164
rect 970 11088 980 11154
rect 1490 11088 1500 11154
rect 970 11078 1500 11088
rect 342 11058 868 11068
rect 342 10992 352 11058
rect 858 10992 868 11058
rect 342 10982 868 10992
rect 970 10962 1500 10972
rect 970 10896 980 10962
rect 1490 10896 1500 10962
rect 970 10886 1500 10896
rect 342 10866 868 10876
rect 342 10800 352 10866
rect 858 10800 868 10866
rect 342 10790 868 10800
rect 970 10770 1500 10780
rect 970 10704 980 10770
rect 1490 10704 1500 10770
rect 970 10694 1500 10704
rect 342 10674 868 10684
rect 342 10608 352 10674
rect 858 10608 868 10674
rect 342 10598 868 10608
rect 970 10578 1500 10588
rect 970 10512 980 10578
rect 1490 10512 1500 10578
rect 970 10502 1500 10512
rect 342 10482 868 10492
rect 342 10416 352 10482
rect 858 10416 868 10482
rect 342 10406 868 10416
rect 970 10386 1500 10396
rect 970 10320 980 10386
rect 1490 10320 1500 10386
rect 970 10310 1500 10320
rect 342 10290 868 10300
rect 342 10224 352 10290
rect 858 10224 868 10290
rect 342 10214 868 10224
rect 970 10194 1500 10204
rect 970 10128 980 10194
rect 1490 10128 1500 10194
rect 970 10118 1500 10128
rect 342 10098 868 10108
rect 342 10032 352 10098
rect 858 10032 868 10098
rect 342 10022 868 10032
rect 970 10002 1500 10012
rect 970 9936 980 10002
rect 1490 9936 1500 10002
rect 970 9926 1500 9936
rect 342 9906 868 9916
rect 342 9840 352 9906
rect 858 9840 868 9906
rect 342 9830 868 9840
rect 970 9810 1500 9820
rect 970 9744 980 9810
rect 1490 9744 1500 9810
rect 970 9734 1500 9744
rect 342 9714 868 9724
rect 342 9648 352 9714
rect 858 9648 868 9714
rect 342 9638 868 9648
rect 970 9618 1500 9628
rect 970 9552 980 9618
rect 1490 9552 1500 9618
rect 970 9542 1500 9552
rect 342 9522 868 9532
rect 342 9456 352 9522
rect 858 9456 868 9522
rect 342 9446 868 9456
rect 970 9426 1500 9436
rect 970 9360 980 9426
rect 1490 9360 1500 9426
rect 970 9350 1500 9360
rect 342 9330 868 9340
rect 342 9264 352 9330
rect 858 9264 868 9330
rect 342 9254 868 9264
rect 970 9234 1500 9244
rect 970 9168 980 9234
rect 1490 9168 1500 9234
rect 970 9158 1500 9168
rect 342 9138 868 9148
rect 342 9072 352 9138
rect 858 9072 868 9138
rect 342 9062 868 9072
rect 970 9042 1500 9052
rect 970 8976 980 9042
rect 1490 8976 1500 9042
rect 970 8966 1500 8976
rect 342 8946 868 8956
rect 342 8880 352 8946
rect 858 8880 868 8946
rect 342 8870 868 8880
rect 970 8850 1500 8860
rect 970 8784 980 8850
rect 1490 8784 1500 8850
rect 970 8774 1500 8784
rect 342 8754 868 8764
rect 342 8688 352 8754
rect 858 8688 868 8754
rect 342 8678 868 8688
rect 970 8658 1500 8668
rect 970 8592 980 8658
rect 1490 8592 1500 8658
rect 970 8582 1500 8592
rect 342 8562 868 8572
rect 342 8496 352 8562
rect 858 8496 868 8562
rect 342 8486 868 8496
rect 970 8466 1500 8476
rect 970 8400 980 8466
rect 1490 8400 1500 8466
rect 970 8390 1500 8400
rect 342 8370 868 8380
rect 342 8304 352 8370
rect 858 8304 868 8370
rect 342 8294 868 8304
rect 970 8274 1500 8284
rect 970 8208 980 8274
rect 1490 8208 1500 8274
rect 970 8198 1500 8208
rect 342 8178 868 8188
rect 342 8112 352 8178
rect 858 8112 868 8178
rect 342 8102 868 8112
rect 970 8082 1500 8092
rect 970 8016 980 8082
rect 1490 8016 1500 8082
rect 970 8006 1500 8016
rect 342 7986 868 7996
rect 342 7920 352 7986
rect 858 7920 868 7986
rect 342 7910 868 7920
rect 970 7890 1500 7900
rect 970 7824 980 7890
rect 1490 7824 1500 7890
rect 970 7814 1500 7824
rect 342 7794 868 7804
rect 342 7728 352 7794
rect 858 7728 868 7794
rect 342 7718 868 7728
rect 970 7698 1500 7708
rect 970 7632 980 7698
rect 1490 7632 1500 7698
rect 970 7622 1500 7632
rect 342 7602 868 7612
rect 342 7536 352 7602
rect 858 7536 868 7602
rect 342 7526 868 7536
rect 970 7506 1500 7516
rect 970 7440 980 7506
rect 1490 7440 1500 7506
rect 970 7430 1500 7440
rect 342 7410 868 7420
rect 342 7344 352 7410
rect 858 7344 868 7410
rect 342 7334 868 7344
rect 970 7314 1500 7324
rect 970 7248 980 7314
rect 1490 7248 1500 7314
rect 970 7238 1500 7248
rect 342 7218 868 7228
rect 342 7152 352 7218
rect 858 7152 868 7218
rect 342 7142 868 7152
rect 970 7122 1500 7132
rect 970 7056 980 7122
rect 1490 7056 1500 7122
rect 970 7046 1500 7056
rect 342 7026 868 7036
rect 342 6960 352 7026
rect 858 6960 868 7026
rect 342 6950 868 6960
rect 970 6930 1500 6940
rect 970 6864 980 6930
rect 1490 6864 1500 6930
rect 970 6854 1500 6864
rect 342 6834 868 6844
rect 342 6768 352 6834
rect 858 6768 868 6834
rect 342 6758 868 6768
rect 970 6738 1500 6748
rect 970 6672 980 6738
rect 1490 6672 1500 6738
rect 970 6662 1500 6672
rect 342 6642 868 6652
rect 342 6576 352 6642
rect 858 6576 868 6642
rect 342 6566 868 6576
rect 970 6546 1500 6556
rect 970 6480 980 6546
rect 1490 6480 1500 6546
rect 970 6470 1500 6480
rect 342 6450 868 6460
rect 342 6384 352 6450
rect 858 6384 868 6450
rect 342 6374 868 6384
rect 970 6354 1500 6364
rect 970 6288 980 6354
rect 1490 6288 1500 6354
rect 970 6278 1500 6288
rect 342 6258 868 6268
rect 342 6192 352 6258
rect 858 6192 868 6258
rect 342 6182 868 6192
rect 970 6162 1500 6172
rect 970 6096 980 6162
rect 1490 6096 1500 6162
rect 970 6086 1500 6096
rect 342 6066 868 6076
rect 342 6000 352 6066
rect 858 6000 868 6066
rect 342 5990 868 6000
rect 970 5970 1500 5980
rect 970 5904 980 5970
rect 1490 5904 1500 5970
rect 970 5894 1500 5904
rect 342 5874 868 5884
rect 342 5808 352 5874
rect 858 5808 868 5874
rect 342 5798 868 5808
rect 970 5778 1500 5788
rect 970 5712 980 5778
rect 1490 5712 1500 5778
rect 970 5702 1500 5712
rect 342 5682 868 5692
rect 342 5616 352 5682
rect 858 5616 868 5682
rect 342 5606 868 5616
rect 970 5586 1500 5596
rect 970 5520 980 5586
rect 1490 5520 1500 5586
rect 970 5510 1500 5520
rect 342 5490 868 5500
rect 342 5424 352 5490
rect 858 5424 868 5490
rect 342 5414 868 5424
rect 970 5394 1500 5404
rect 970 5328 980 5394
rect 1490 5328 1500 5394
rect 970 5318 1500 5328
rect 342 5298 868 5308
rect 342 5232 352 5298
rect 858 5232 868 5298
rect 342 5222 868 5232
rect 970 5202 1500 5212
rect 970 5136 980 5202
rect 1490 5136 1500 5202
rect 970 5126 1500 5136
rect 342 5106 868 5116
rect 342 5040 352 5106
rect 858 5040 868 5106
rect 342 5030 868 5040
rect 970 5010 1500 5020
rect 970 4944 980 5010
rect 1490 4944 1500 5010
rect 970 4934 1500 4944
rect 342 4914 868 4924
rect 342 4848 352 4914
rect 858 4848 868 4914
rect 342 4838 868 4848
rect 970 4818 1500 4828
rect 970 4752 980 4818
rect 1490 4752 1500 4818
rect 970 4742 1500 4752
rect 342 4722 868 4732
rect 342 4656 352 4722
rect 858 4656 868 4722
rect 342 4646 868 4656
rect 970 4626 1500 4636
rect 970 4560 980 4626
rect 1490 4560 1500 4626
rect 970 4550 1500 4560
rect 342 4530 868 4540
rect 342 4464 352 4530
rect 858 4464 868 4530
rect 342 4454 868 4464
rect 970 4434 1500 4444
rect 970 4368 980 4434
rect 1490 4368 1500 4434
rect 970 4358 1500 4368
rect 342 4338 868 4348
rect 342 4272 352 4338
rect 858 4272 868 4338
rect 342 4262 868 4272
rect 970 4242 1500 4252
rect 970 4176 980 4242
rect 1490 4176 1500 4242
rect 970 4166 1500 4176
rect 342 4146 868 4156
rect 342 4080 352 4146
rect 858 4080 868 4146
rect 342 4070 868 4080
rect 970 4050 1500 4060
rect 970 3984 980 4050
rect 1490 3984 1500 4050
rect 970 3974 1500 3984
rect 342 3954 868 3964
rect 342 3888 352 3954
rect 858 3888 868 3954
rect 342 3878 868 3888
rect 970 3858 1500 3868
rect 970 3792 980 3858
rect 1490 3792 1500 3858
rect 970 3782 1500 3792
rect 342 3762 868 3772
rect 342 3696 352 3762
rect 858 3696 868 3762
rect 342 3686 868 3696
rect 970 3666 1500 3676
rect 970 3600 980 3666
rect 1490 3600 1500 3666
rect 970 3590 1500 3600
rect 342 3570 868 3580
rect 342 3504 352 3570
rect 858 3504 868 3570
rect 342 3494 868 3504
rect 970 3474 1500 3484
rect 970 3408 980 3474
rect 1490 3408 1500 3474
rect 970 3398 1500 3408
rect 342 3378 868 3388
rect 342 3312 352 3378
rect 858 3312 868 3378
rect 342 3302 868 3312
rect 970 3282 1500 3292
rect 970 3216 980 3282
rect 1490 3216 1500 3282
rect 970 3206 1500 3216
rect 342 3186 868 3196
rect 342 3120 352 3186
rect 858 3120 868 3186
rect 342 3110 868 3120
rect 970 3090 1500 3100
rect 970 3024 980 3090
rect 1490 3024 1500 3090
rect 970 3014 1500 3024
rect 342 2994 868 3004
rect 342 2928 352 2994
rect 858 2928 868 2994
rect 342 2918 868 2928
rect 970 2898 1500 2908
rect 970 2832 980 2898
rect 1490 2832 1500 2898
rect 970 2822 1500 2832
rect 342 2802 868 2812
rect 342 2736 352 2802
rect 858 2736 868 2802
rect 342 2726 868 2736
rect 970 2706 1500 2716
rect 970 2640 980 2706
rect 1490 2640 1500 2706
rect 970 2630 1500 2640
rect 342 2610 868 2620
rect 342 2544 352 2610
rect 858 2544 868 2610
rect 342 2534 868 2544
rect 970 2514 1500 2524
rect 970 2448 980 2514
rect 1490 2448 1500 2514
rect 970 2438 1500 2448
rect 342 2418 868 2428
rect 342 2352 352 2418
rect 858 2352 868 2418
rect 342 2342 868 2352
rect 970 2322 1500 2332
rect 970 2256 980 2322
rect 1490 2256 1500 2322
rect 970 2246 1500 2256
rect 342 2226 868 2236
rect 342 2160 352 2226
rect 858 2160 868 2226
rect 342 2150 868 2160
rect 970 2130 1500 2140
rect 970 2064 980 2130
rect 1490 2064 1500 2130
rect 970 2054 1500 2064
rect 342 2034 868 2044
rect 342 1968 352 2034
rect 858 1968 868 2034
rect 342 1958 868 1968
rect 970 1938 1500 1948
rect 970 1872 980 1938
rect 1490 1872 1500 1938
rect 970 1862 1500 1872
rect 342 1842 868 1852
rect 342 1776 352 1842
rect 858 1776 868 1842
rect 342 1766 868 1776
rect 970 1746 1500 1756
rect 970 1680 980 1746
rect 1490 1680 1500 1746
rect 970 1670 1500 1680
rect 342 1650 868 1660
rect 342 1584 352 1650
rect 858 1584 868 1650
rect 342 1574 868 1584
rect 970 1554 1500 1564
rect 970 1488 980 1554
rect 1490 1488 1500 1554
rect 970 1478 1500 1488
rect 342 1458 868 1468
rect 342 1392 352 1458
rect 858 1392 868 1458
rect 342 1382 868 1392
rect 970 1362 1500 1372
rect 970 1296 980 1362
rect 1490 1296 1500 1362
rect 970 1286 1500 1296
rect 342 1266 868 1276
rect 342 1200 352 1266
rect 858 1200 868 1266
rect 342 1190 868 1200
rect 970 1170 1500 1180
rect 970 1104 980 1170
rect 1490 1104 1500 1170
rect 970 1094 1500 1104
rect 342 1074 868 1084
rect 342 1008 352 1074
rect 858 1008 868 1074
rect 342 998 868 1008
rect 970 978 1500 988
rect 970 912 980 978
rect 1490 912 1500 978
rect 970 902 1500 912
rect 342 882 868 892
rect 342 816 352 882
rect 858 816 868 882
rect 342 806 868 816
rect 970 786 1500 796
rect 970 720 980 786
rect 1490 720 1500 786
rect 970 710 1500 720
rect 342 690 868 700
rect 342 624 352 690
rect 858 624 868 690
rect 342 614 868 624
<< via2 >>
rect 132 22222 1706 22286
rect 352 21868 858 21934
rect 352 21744 858 21810
rect 980 21648 1490 21714
rect 352 21552 858 21618
rect 980 21456 1490 21522
rect 352 21360 858 21426
rect 980 21264 1490 21330
rect 352 21168 858 21234
rect 980 21072 1490 21138
rect 352 20976 858 21042
rect 980 20880 1490 20946
rect 352 20784 858 20850
rect 980 20688 1490 20754
rect 352 20592 858 20658
rect 980 20496 1490 20562
rect 352 20400 858 20466
rect 980 20304 1490 20370
rect 352 20208 858 20274
rect 980 20112 1490 20178
rect 352 20016 858 20082
rect 980 19920 1490 19986
rect 352 19824 858 19890
rect 980 19728 1490 19794
rect 352 19632 858 19698
rect 980 19536 1490 19602
rect 352 19440 858 19506
rect 980 19344 1490 19410
rect 352 19248 858 19314
rect 980 19152 1490 19218
rect 352 19056 858 19122
rect 980 18960 1490 19026
rect 352 18864 858 18930
rect 980 18768 1490 18834
rect 352 18672 858 18738
rect 980 18576 1490 18642
rect 352 18480 858 18546
rect 980 18384 1490 18450
rect 352 18288 858 18354
rect 980 18192 1490 18258
rect 352 18096 858 18162
rect 980 18000 1490 18066
rect 352 17904 858 17970
rect 980 17808 1490 17874
rect 352 17712 858 17778
rect 980 17616 1490 17682
rect 352 17520 858 17586
rect 980 17424 1490 17490
rect 352 17328 858 17394
rect 980 17232 1490 17298
rect 352 17136 858 17202
rect 980 17040 1490 17106
rect 352 16944 858 17010
rect 980 16848 1490 16914
rect 352 16752 858 16818
rect 980 16656 1490 16722
rect 352 16560 858 16626
rect 980 16464 1490 16530
rect 352 16368 858 16434
rect 980 16272 1490 16338
rect 352 16176 858 16242
rect 980 16080 1490 16146
rect 352 15984 858 16050
rect 980 15888 1490 15954
rect 352 15792 858 15858
rect 980 15696 1490 15762
rect 352 15600 858 15666
rect 980 15504 1490 15570
rect 352 15408 858 15474
rect 980 15312 1490 15378
rect 352 15216 858 15282
rect 980 15120 1490 15186
rect 352 15024 858 15090
rect 980 14928 1490 14994
rect 352 14832 858 14898
rect 980 14736 1490 14802
rect 352 14640 858 14706
rect 980 14544 1490 14610
rect 352 14448 858 14514
rect 980 14352 1490 14418
rect 352 14256 858 14322
rect 980 14160 1490 14226
rect 352 14064 858 14130
rect 980 13968 1490 14034
rect 352 13872 858 13938
rect 980 13776 1490 13842
rect 352 13680 858 13746
rect 980 13584 1490 13650
rect 352 13488 858 13554
rect 980 13392 1490 13458
rect 352 13296 858 13362
rect 980 13200 1490 13266
rect 352 13104 858 13170
rect 980 13008 1490 13074
rect 352 12912 858 12978
rect 980 12816 1490 12882
rect 352 12720 858 12786
rect 980 12624 1490 12690
rect 352 12528 858 12594
rect 980 12432 1490 12498
rect 352 12336 858 12402
rect 980 12240 1490 12306
rect 352 12144 858 12210
rect 980 12048 1490 12114
rect 352 11952 858 12018
rect 980 11856 1490 11922
rect 352 11760 858 11826
rect 980 11664 1490 11730
rect 352 11568 858 11634
rect 980 11472 1490 11538
rect 352 11376 858 11442
rect 980 11280 1490 11346
rect 352 11184 858 11250
rect 980 11088 1490 11154
rect 352 10992 858 11058
rect 980 10896 1490 10962
rect 352 10800 858 10866
rect 980 10704 1490 10770
rect 352 10608 858 10674
rect 980 10512 1490 10578
rect 352 10416 858 10482
rect 980 10320 1490 10386
rect 352 10224 858 10290
rect 980 10128 1490 10194
rect 352 10032 858 10098
rect 980 9936 1490 10002
rect 352 9840 858 9906
rect 980 9744 1490 9810
rect 352 9648 858 9714
rect 980 9552 1490 9618
rect 352 9456 858 9522
rect 980 9360 1490 9426
rect 352 9264 858 9330
rect 980 9168 1490 9234
rect 352 9072 858 9138
rect 980 8976 1490 9042
rect 352 8880 858 8946
rect 980 8784 1490 8850
rect 352 8688 858 8754
rect 980 8592 1490 8658
rect 352 8496 858 8562
rect 980 8400 1490 8466
rect 352 8304 858 8370
rect 980 8208 1490 8274
rect 352 8112 858 8178
rect 980 8016 1490 8082
rect 352 7920 858 7986
rect 980 7824 1490 7890
rect 352 7728 858 7794
rect 980 7632 1490 7698
rect 352 7536 858 7602
rect 980 7440 1490 7506
rect 352 7344 858 7410
rect 980 7248 1490 7314
rect 352 7152 858 7218
rect 980 7056 1490 7122
rect 352 6960 858 7026
rect 980 6864 1490 6930
rect 352 6768 858 6834
rect 980 6672 1490 6738
rect 352 6576 858 6642
rect 980 6480 1490 6546
rect 352 6384 858 6450
rect 980 6288 1490 6354
rect 352 6192 858 6258
rect 980 6096 1490 6162
rect 352 6000 858 6066
rect 980 5904 1490 5970
rect 352 5808 858 5874
rect 980 5712 1490 5778
rect 352 5616 858 5682
rect 980 5520 1490 5586
rect 352 5424 858 5490
rect 980 5328 1490 5394
rect 352 5232 858 5298
rect 980 5136 1490 5202
rect 352 5040 858 5106
rect 980 4944 1490 5010
rect 352 4848 858 4914
rect 980 4752 1490 4818
rect 352 4656 858 4722
rect 980 4560 1490 4626
rect 352 4464 858 4530
rect 980 4368 1490 4434
rect 352 4272 858 4338
rect 980 4176 1490 4242
rect 352 4080 858 4146
rect 980 3984 1490 4050
rect 352 3888 858 3954
rect 980 3792 1490 3858
rect 352 3696 858 3762
rect 980 3600 1490 3666
rect 352 3504 858 3570
rect 980 3408 1490 3474
rect 352 3312 858 3378
rect 980 3216 1490 3282
rect 352 3120 858 3186
rect 980 3024 1490 3090
rect 352 2928 858 2994
rect 980 2832 1490 2898
rect 352 2736 858 2802
rect 980 2640 1490 2706
rect 352 2544 858 2610
rect 980 2448 1490 2514
rect 352 2352 858 2418
rect 980 2256 1490 2322
rect 352 2160 858 2226
rect 980 2064 1490 2130
rect 352 1968 858 2034
rect 980 1872 1490 1938
rect 352 1776 858 1842
rect 980 1680 1490 1746
rect 352 1584 858 1650
rect 980 1488 1490 1554
rect 352 1392 858 1458
rect 980 1296 1490 1362
rect 352 1200 858 1266
rect 980 1104 1490 1170
rect 352 1008 858 1074
rect 980 912 1490 978
rect 352 816 858 882
rect 980 720 1490 786
rect 352 624 858 690
<< metal3 >>
rect 122 22286 1716 22291
rect 122 22222 132 22286
rect 1706 22222 1716 22286
rect 122 22217 1716 22222
rect 344 21934 868 21944
rect 344 21868 352 21934
rect 858 21868 868 21934
rect 344 21820 868 21868
rect 342 21810 868 21820
rect 342 21744 352 21810
rect 858 21744 868 21810
rect 342 21734 868 21744
rect 970 21714 1500 21724
rect 970 21648 980 21714
rect 1490 21648 1500 21714
rect 970 21638 1500 21648
rect 342 21618 868 21628
rect 342 21552 352 21618
rect 858 21552 868 21618
rect 342 21542 868 21552
rect 970 21522 1500 21532
rect 970 21456 980 21522
rect 1490 21456 1500 21522
rect 970 21446 1500 21456
rect 342 21426 868 21436
rect 342 21360 352 21426
rect 858 21360 868 21426
rect 342 21350 868 21360
rect 970 21330 1500 21340
rect 970 21264 980 21330
rect 1490 21264 1500 21330
rect 970 21254 1500 21264
rect 342 21234 868 21244
rect 342 21168 352 21234
rect 858 21168 868 21234
rect 342 21158 868 21168
rect 970 21138 1500 21148
rect 970 21072 980 21138
rect 1490 21072 1500 21138
rect 970 21062 1500 21072
rect 342 21042 868 21052
rect 342 20976 352 21042
rect 858 20976 868 21042
rect 342 20966 868 20976
rect 970 20946 1500 20956
rect 970 20880 980 20946
rect 1490 20880 1500 20946
rect 970 20870 1500 20880
rect 342 20850 868 20860
rect 342 20784 352 20850
rect 858 20784 868 20850
rect 342 20774 868 20784
rect 970 20754 1500 20764
rect 970 20688 980 20754
rect 1490 20688 1500 20754
rect 970 20678 1500 20688
rect 342 20658 868 20668
rect 342 20592 352 20658
rect 858 20592 868 20658
rect 342 20582 868 20592
rect 970 20562 1500 20572
rect 970 20496 980 20562
rect 1490 20496 1500 20562
rect 970 20486 1500 20496
rect 342 20466 868 20476
rect 342 20400 352 20466
rect 858 20400 868 20466
rect 342 20390 868 20400
rect 970 20370 1500 20380
rect 970 20304 980 20370
rect 1490 20304 1500 20370
rect 970 20294 1500 20304
rect 342 20274 868 20284
rect 342 20208 352 20274
rect 858 20208 868 20274
rect 342 20198 868 20208
rect 970 20178 1500 20188
rect 970 20112 980 20178
rect 1490 20112 1500 20178
rect 970 20102 1500 20112
rect 342 20082 868 20092
rect 342 20016 352 20082
rect 858 20016 868 20082
rect 342 20006 868 20016
rect 970 19986 1500 19996
rect 970 19920 980 19986
rect 1490 19920 1500 19986
rect 970 19910 1500 19920
rect 342 19890 868 19900
rect 342 19824 352 19890
rect 858 19824 868 19890
rect 342 19814 868 19824
rect 970 19794 1500 19804
rect 970 19728 980 19794
rect 1490 19728 1500 19794
rect 970 19718 1500 19728
rect 342 19698 868 19708
rect 342 19632 352 19698
rect 858 19632 868 19698
rect 342 19622 868 19632
rect 970 19602 1500 19612
rect 970 19536 980 19602
rect 1490 19536 1500 19602
rect 970 19526 1500 19536
rect 342 19506 868 19516
rect 342 19440 352 19506
rect 858 19440 868 19506
rect 342 19430 868 19440
rect 970 19410 1500 19420
rect 970 19344 980 19410
rect 1490 19344 1500 19410
rect 970 19334 1500 19344
rect 342 19314 868 19324
rect 342 19248 352 19314
rect 858 19248 868 19314
rect 342 19238 868 19248
rect 970 19218 1500 19228
rect 970 19152 980 19218
rect 1490 19152 1500 19218
rect 970 19142 1500 19152
rect 342 19122 868 19132
rect 342 19056 352 19122
rect 858 19056 868 19122
rect 342 19046 868 19056
rect 970 19026 1500 19036
rect 970 18960 980 19026
rect 1490 18960 1500 19026
rect 970 18950 1500 18960
rect 342 18930 868 18940
rect 342 18864 352 18930
rect 858 18864 868 18930
rect 342 18854 868 18864
rect 970 18834 1500 18844
rect 970 18768 980 18834
rect 1490 18768 1500 18834
rect 970 18758 1500 18768
rect 342 18738 868 18748
rect 342 18672 352 18738
rect 858 18672 868 18738
rect 342 18662 868 18672
rect 970 18642 1500 18652
rect 970 18576 980 18642
rect 1490 18576 1500 18642
rect 970 18566 1500 18576
rect 342 18546 868 18556
rect 342 18480 352 18546
rect 858 18480 868 18546
rect 342 18470 868 18480
rect 970 18450 1500 18460
rect 970 18384 980 18450
rect 1490 18384 1500 18450
rect 970 18374 1500 18384
rect 342 18354 868 18364
rect 342 18288 352 18354
rect 858 18288 868 18354
rect 342 18278 868 18288
rect 970 18258 1500 18268
rect 970 18192 980 18258
rect 1490 18192 1500 18258
rect 970 18182 1500 18192
rect 342 18162 868 18172
rect 342 18096 352 18162
rect 858 18096 868 18162
rect 342 18086 868 18096
rect 970 18066 1500 18076
rect 970 18000 980 18066
rect 1490 18000 1500 18066
rect 970 17990 1500 18000
rect 342 17970 868 17980
rect 342 17904 352 17970
rect 858 17904 868 17970
rect 342 17894 868 17904
rect 970 17874 1500 17884
rect 970 17808 980 17874
rect 1490 17808 1500 17874
rect 970 17798 1500 17808
rect 342 17778 868 17788
rect 342 17712 352 17778
rect 858 17712 868 17778
rect 342 17702 868 17712
rect 970 17682 1500 17692
rect 970 17616 980 17682
rect 1490 17616 1500 17682
rect 970 17606 1500 17616
rect 342 17586 868 17596
rect 342 17520 352 17586
rect 858 17520 868 17586
rect 342 17510 868 17520
rect 970 17490 1500 17500
rect 970 17424 980 17490
rect 1490 17424 1500 17490
rect 970 17414 1500 17424
rect 342 17394 868 17404
rect 342 17328 352 17394
rect 858 17328 868 17394
rect 342 17318 868 17328
rect 970 17298 1500 17308
rect 970 17232 980 17298
rect 1490 17232 1500 17298
rect 970 17222 1500 17232
rect 342 17202 868 17212
rect 342 17136 352 17202
rect 858 17136 868 17202
rect 342 17126 868 17136
rect 970 17106 1500 17116
rect 970 17040 980 17106
rect 1490 17040 1500 17106
rect 970 17030 1500 17040
rect 342 17010 868 17020
rect 342 16944 352 17010
rect 858 16944 868 17010
rect 342 16934 868 16944
rect 970 16914 1500 16924
rect 970 16848 980 16914
rect 1490 16848 1500 16914
rect 970 16838 1500 16848
rect 342 16818 868 16828
rect 342 16752 352 16818
rect 858 16752 868 16818
rect 342 16742 868 16752
rect 970 16722 1500 16732
rect 970 16656 980 16722
rect 1490 16656 1500 16722
rect 970 16646 1500 16656
rect 342 16626 868 16636
rect 342 16560 352 16626
rect 858 16560 868 16626
rect 342 16550 868 16560
rect 970 16530 1500 16540
rect 970 16464 980 16530
rect 1490 16464 1500 16530
rect 970 16454 1500 16464
rect 342 16434 868 16444
rect 342 16368 352 16434
rect 858 16368 868 16434
rect 342 16358 868 16368
rect 970 16338 1500 16348
rect 970 16272 980 16338
rect 1490 16272 1500 16338
rect 970 16262 1500 16272
rect 342 16242 868 16252
rect 342 16176 352 16242
rect 858 16176 868 16242
rect 342 16166 868 16176
rect 970 16146 1500 16156
rect 970 16080 980 16146
rect 1490 16080 1500 16146
rect 970 16070 1500 16080
rect 342 16050 868 16060
rect 342 15984 352 16050
rect 858 15984 868 16050
rect 342 15974 868 15984
rect 970 15954 1500 15964
rect 970 15888 980 15954
rect 1490 15888 1500 15954
rect 970 15878 1500 15888
rect 342 15858 868 15868
rect 342 15792 352 15858
rect 858 15792 868 15858
rect 342 15782 868 15792
rect 970 15762 1500 15772
rect 970 15696 980 15762
rect 1490 15696 1500 15762
rect 970 15686 1500 15696
rect 342 15666 868 15676
rect 342 15600 352 15666
rect 858 15600 868 15666
rect 342 15590 868 15600
rect 970 15570 1500 15580
rect 970 15504 980 15570
rect 1490 15504 1500 15570
rect 970 15494 1500 15504
rect 342 15474 868 15484
rect 342 15408 352 15474
rect 858 15408 868 15474
rect 342 15398 868 15408
rect 970 15378 1500 15388
rect 970 15312 980 15378
rect 1490 15312 1500 15378
rect 970 15302 1500 15312
rect 342 15282 868 15292
rect 342 15216 352 15282
rect 858 15216 868 15282
rect 342 15206 868 15216
rect 970 15186 1500 15196
rect 970 15120 980 15186
rect 1490 15120 1500 15186
rect 970 15110 1500 15120
rect 342 15090 868 15100
rect 342 15024 352 15090
rect 858 15024 868 15090
rect 342 15014 868 15024
rect 970 14994 1500 15004
rect 970 14928 980 14994
rect 1490 14928 1500 14994
rect 970 14918 1500 14928
rect 342 14898 868 14908
rect 342 14832 352 14898
rect 858 14832 868 14898
rect 342 14822 868 14832
rect 970 14802 1500 14812
rect 970 14736 980 14802
rect 1490 14736 1500 14802
rect 970 14726 1500 14736
rect 342 14706 868 14716
rect 342 14640 352 14706
rect 858 14640 868 14706
rect 342 14630 868 14640
rect 970 14610 1500 14620
rect 970 14544 980 14610
rect 1490 14544 1500 14610
rect 970 14534 1500 14544
rect 342 14514 868 14524
rect 342 14448 352 14514
rect 858 14448 868 14514
rect 342 14438 868 14448
rect 970 14418 1500 14428
rect 970 14352 980 14418
rect 1490 14352 1500 14418
rect 970 14342 1500 14352
rect 342 14322 868 14332
rect 342 14256 352 14322
rect 858 14256 868 14322
rect 342 14246 868 14256
rect 970 14226 1500 14236
rect 970 14160 980 14226
rect 1490 14160 1500 14226
rect 970 14150 1500 14160
rect 342 14130 868 14140
rect 342 14064 352 14130
rect 858 14064 868 14130
rect 342 14054 868 14064
rect 970 14034 1500 14044
rect 970 13968 980 14034
rect 1490 13968 1500 14034
rect 970 13958 1500 13968
rect 342 13938 868 13948
rect 342 13872 352 13938
rect 858 13872 868 13938
rect 342 13862 868 13872
rect 970 13842 1500 13852
rect 970 13776 980 13842
rect 1490 13776 1500 13842
rect 970 13766 1500 13776
rect 342 13746 868 13756
rect 342 13680 352 13746
rect 858 13680 868 13746
rect 342 13670 868 13680
rect 970 13650 1500 13660
rect 970 13584 980 13650
rect 1490 13584 1500 13650
rect 970 13574 1500 13584
rect 342 13554 868 13564
rect 342 13488 352 13554
rect 858 13488 868 13554
rect 342 13478 868 13488
rect 970 13458 1500 13468
rect 970 13392 980 13458
rect 1490 13392 1500 13458
rect 970 13382 1500 13392
rect 342 13362 868 13372
rect 342 13296 352 13362
rect 858 13296 868 13362
rect 342 13286 868 13296
rect 970 13266 1500 13276
rect 970 13200 980 13266
rect 1490 13200 1500 13266
rect 970 13190 1500 13200
rect 342 13170 868 13180
rect 342 13104 352 13170
rect 858 13104 868 13170
rect 342 13094 868 13104
rect 970 13074 1500 13084
rect 970 13008 980 13074
rect 1490 13008 1500 13074
rect 970 12998 1500 13008
rect 342 12978 868 12988
rect 342 12912 352 12978
rect 858 12912 868 12978
rect 342 12902 868 12912
rect 970 12882 1500 12892
rect 970 12816 980 12882
rect 1490 12816 1500 12882
rect 970 12806 1500 12816
rect 342 12786 868 12796
rect 342 12720 352 12786
rect 858 12720 868 12786
rect 342 12710 868 12720
rect 970 12690 1500 12700
rect 970 12624 980 12690
rect 1490 12624 1500 12690
rect 970 12614 1500 12624
rect 342 12594 868 12604
rect 342 12528 352 12594
rect 858 12528 868 12594
rect 342 12518 868 12528
rect 970 12498 1500 12508
rect 970 12432 980 12498
rect 1490 12432 1500 12498
rect 970 12422 1500 12432
rect 342 12402 868 12412
rect 342 12336 352 12402
rect 858 12336 868 12402
rect 342 12326 868 12336
rect 970 12306 1500 12316
rect 970 12240 980 12306
rect 1490 12240 1500 12306
rect 970 12230 1500 12240
rect 342 12210 868 12220
rect 342 12144 352 12210
rect 858 12144 868 12210
rect 342 12134 868 12144
rect 970 12114 1500 12124
rect 970 12048 980 12114
rect 1490 12048 1500 12114
rect 970 12038 1500 12048
rect 342 12018 868 12028
rect 342 11952 352 12018
rect 858 11952 868 12018
rect 342 11942 868 11952
rect 970 11922 1500 11932
rect 970 11856 980 11922
rect 1490 11856 1500 11922
rect 970 11846 1500 11856
rect 342 11826 868 11836
rect 342 11760 352 11826
rect 858 11760 868 11826
rect 342 11750 868 11760
rect 970 11730 1500 11740
rect 970 11664 980 11730
rect 1490 11664 1500 11730
rect 970 11654 1500 11664
rect 342 11634 868 11644
rect 342 11568 352 11634
rect 858 11568 868 11634
rect 342 11558 868 11568
rect 970 11538 1500 11548
rect 970 11472 980 11538
rect 1490 11472 1500 11538
rect 970 11462 1500 11472
rect 342 11442 868 11452
rect 342 11376 352 11442
rect 858 11376 868 11442
rect 342 11366 868 11376
rect 970 11346 1500 11356
rect 970 11280 980 11346
rect 1490 11280 1500 11346
rect 970 11270 1500 11280
rect 342 11250 868 11260
rect 342 11184 352 11250
rect 858 11184 868 11250
rect 342 11174 868 11184
rect 970 11154 1500 11164
rect 970 11088 980 11154
rect 1490 11088 1500 11154
rect 970 11078 1500 11088
rect 342 11058 868 11068
rect 342 10992 352 11058
rect 858 10992 868 11058
rect 342 10982 868 10992
rect 970 10962 1500 10972
rect 970 10896 980 10962
rect 1490 10896 1500 10962
rect 970 10886 1500 10896
rect 342 10866 868 10876
rect 342 10800 352 10866
rect 858 10800 868 10866
rect 342 10790 868 10800
rect 970 10770 1500 10780
rect 970 10704 980 10770
rect 1490 10704 1500 10770
rect 970 10694 1500 10704
rect 342 10674 868 10684
rect 342 10608 352 10674
rect 858 10608 868 10674
rect 342 10598 868 10608
rect 970 10578 1500 10588
rect 970 10512 980 10578
rect 1490 10512 1500 10578
rect 970 10502 1500 10512
rect 342 10482 868 10492
rect 342 10416 352 10482
rect 858 10416 868 10482
rect 342 10406 868 10416
rect 970 10386 1500 10396
rect 970 10320 980 10386
rect 1490 10320 1500 10386
rect 970 10310 1500 10320
rect 342 10290 868 10300
rect 342 10224 352 10290
rect 858 10224 868 10290
rect 342 10214 868 10224
rect 970 10194 1500 10204
rect 970 10128 980 10194
rect 1490 10128 1500 10194
rect 970 10118 1500 10128
rect 342 10098 868 10108
rect 342 10032 352 10098
rect 858 10032 868 10098
rect 342 10022 868 10032
rect 970 10002 1500 10012
rect 970 9936 980 10002
rect 1490 9936 1500 10002
rect 970 9926 1500 9936
rect 342 9906 868 9916
rect 342 9840 352 9906
rect 858 9840 868 9906
rect 342 9830 868 9840
rect 970 9810 1500 9820
rect 970 9744 980 9810
rect 1490 9744 1500 9810
rect 970 9734 1500 9744
rect 342 9714 868 9724
rect 342 9648 352 9714
rect 858 9648 868 9714
rect 342 9638 868 9648
rect 970 9618 1500 9628
rect 970 9552 980 9618
rect 1490 9552 1500 9618
rect 970 9542 1500 9552
rect 342 9522 868 9532
rect 342 9456 352 9522
rect 858 9456 868 9522
rect 342 9446 868 9456
rect 970 9426 1500 9436
rect 970 9360 980 9426
rect 1490 9360 1500 9426
rect 970 9350 1500 9360
rect 342 9330 868 9340
rect 342 9264 352 9330
rect 858 9264 868 9330
rect 342 9254 868 9264
rect 970 9234 1500 9244
rect 970 9168 980 9234
rect 1490 9168 1500 9234
rect 970 9158 1500 9168
rect 342 9138 868 9148
rect 342 9072 352 9138
rect 858 9072 868 9138
rect 342 9062 868 9072
rect 970 9042 1500 9052
rect 970 8976 980 9042
rect 1490 8976 1500 9042
rect 970 8966 1500 8976
rect 342 8946 868 8956
rect 342 8880 352 8946
rect 858 8880 868 8946
rect 342 8870 868 8880
rect 970 8850 1500 8860
rect 970 8784 980 8850
rect 1490 8784 1500 8850
rect 970 8774 1500 8784
rect 342 8754 868 8764
rect 342 8688 352 8754
rect 858 8688 868 8754
rect 342 8678 868 8688
rect 970 8658 1500 8668
rect 970 8592 980 8658
rect 1490 8592 1500 8658
rect 970 8582 1500 8592
rect 342 8562 868 8572
rect 342 8496 352 8562
rect 858 8496 868 8562
rect 342 8486 868 8496
rect 970 8466 1500 8476
rect 970 8400 980 8466
rect 1490 8400 1500 8466
rect 970 8390 1500 8400
rect 342 8370 868 8380
rect 342 8304 352 8370
rect 858 8304 868 8370
rect 342 8294 868 8304
rect 970 8274 1500 8284
rect 970 8208 980 8274
rect 1490 8208 1500 8274
rect 970 8198 1500 8208
rect 342 8178 868 8188
rect 342 8112 352 8178
rect 858 8112 868 8178
rect 342 8102 868 8112
rect 970 8082 1500 8092
rect 970 8016 980 8082
rect 1490 8016 1500 8082
rect 970 8006 1500 8016
rect 342 7986 868 7996
rect 342 7920 352 7986
rect 858 7920 868 7986
rect 342 7910 868 7920
rect 970 7890 1500 7900
rect 970 7824 980 7890
rect 1490 7824 1500 7890
rect 970 7814 1500 7824
rect 342 7794 868 7804
rect 342 7728 352 7794
rect 858 7728 868 7794
rect 342 7718 868 7728
rect 970 7698 1500 7708
rect 970 7632 980 7698
rect 1490 7632 1500 7698
rect 970 7622 1500 7632
rect 342 7602 868 7612
rect 342 7536 352 7602
rect 858 7536 868 7602
rect 342 7526 868 7536
rect 970 7506 1500 7516
rect 970 7440 980 7506
rect 1490 7440 1500 7506
rect 970 7430 1500 7440
rect 342 7410 868 7420
rect 342 7344 352 7410
rect 858 7344 868 7410
rect 342 7334 868 7344
rect 970 7314 1500 7324
rect 970 7248 980 7314
rect 1490 7248 1500 7314
rect 970 7238 1500 7248
rect 342 7218 868 7228
rect 342 7152 352 7218
rect 858 7152 868 7218
rect 342 7142 868 7152
rect 970 7122 1500 7132
rect 970 7056 980 7122
rect 1490 7056 1500 7122
rect 970 7046 1500 7056
rect 342 7026 868 7036
rect 342 6960 352 7026
rect 858 6960 868 7026
rect 342 6950 868 6960
rect 970 6930 1500 6940
rect 970 6864 980 6930
rect 1490 6864 1500 6930
rect 970 6854 1500 6864
rect 342 6834 868 6844
rect 342 6768 352 6834
rect 858 6768 868 6834
rect 342 6758 868 6768
rect 970 6738 1500 6748
rect 970 6672 980 6738
rect 1490 6672 1500 6738
rect 970 6662 1500 6672
rect 342 6642 868 6652
rect 342 6576 352 6642
rect 858 6576 868 6642
rect 342 6566 868 6576
rect 970 6546 1500 6556
rect 970 6480 980 6546
rect 1490 6480 1500 6546
rect 970 6470 1500 6480
rect 342 6450 868 6460
rect 342 6384 352 6450
rect 858 6384 868 6450
rect 342 6374 868 6384
rect 970 6354 1500 6364
rect 970 6288 980 6354
rect 1490 6288 1500 6354
rect 970 6278 1500 6288
rect 342 6258 868 6268
rect 342 6192 352 6258
rect 858 6192 868 6258
rect 342 6182 868 6192
rect 970 6162 1500 6172
rect 970 6096 980 6162
rect 1490 6096 1500 6162
rect 970 6086 1500 6096
rect 342 6066 868 6076
rect 342 6000 352 6066
rect 858 6000 868 6066
rect 342 5990 868 6000
rect 970 5970 1500 5980
rect 970 5904 980 5970
rect 1490 5904 1500 5970
rect 970 5894 1500 5904
rect 342 5874 868 5884
rect 342 5808 352 5874
rect 858 5808 868 5874
rect 342 5798 868 5808
rect 970 5778 1500 5788
rect 970 5712 980 5778
rect 1490 5712 1500 5778
rect 970 5702 1500 5712
rect 342 5682 868 5692
rect 342 5616 352 5682
rect 858 5616 868 5682
rect 342 5606 868 5616
rect 970 5586 1500 5596
rect 970 5520 980 5586
rect 1490 5520 1500 5586
rect 970 5510 1500 5520
rect 342 5490 868 5500
rect 342 5424 352 5490
rect 858 5424 868 5490
rect 342 5414 868 5424
rect 970 5394 1500 5404
rect 970 5328 980 5394
rect 1490 5328 1500 5394
rect 970 5318 1500 5328
rect 342 5298 868 5308
rect 342 5232 352 5298
rect 858 5232 868 5298
rect 342 5222 868 5232
rect 970 5202 1500 5212
rect 970 5136 980 5202
rect 1490 5136 1500 5202
rect 970 5126 1500 5136
rect 342 5106 868 5116
rect 342 5040 352 5106
rect 858 5040 868 5106
rect 342 5030 868 5040
rect 970 5010 1500 5020
rect 970 4944 980 5010
rect 1490 4944 1500 5010
rect 970 4934 1500 4944
rect 342 4914 868 4924
rect 342 4848 352 4914
rect 858 4848 868 4914
rect 342 4838 868 4848
rect 970 4818 1500 4828
rect 970 4752 980 4818
rect 1490 4752 1500 4818
rect 970 4742 1500 4752
rect 342 4722 868 4732
rect 342 4656 352 4722
rect 858 4656 868 4722
rect 342 4646 868 4656
rect 970 4626 1500 4636
rect 970 4560 980 4626
rect 1490 4560 1500 4626
rect 970 4550 1500 4560
rect 342 4530 868 4540
rect 342 4464 352 4530
rect 858 4464 868 4530
rect 342 4454 868 4464
rect 970 4434 1500 4444
rect 970 4368 980 4434
rect 1490 4368 1500 4434
rect 970 4358 1500 4368
rect 342 4338 868 4348
rect 342 4272 352 4338
rect 858 4272 868 4338
rect 342 4262 868 4272
rect 970 4242 1500 4252
rect 970 4176 980 4242
rect 1490 4176 1500 4242
rect 970 4166 1500 4176
rect 342 4146 868 4156
rect 342 4080 352 4146
rect 858 4080 868 4146
rect 342 4070 868 4080
rect 970 4050 1500 4060
rect 970 3984 980 4050
rect 1490 3984 1500 4050
rect 970 3974 1500 3984
rect 342 3954 868 3964
rect 342 3888 352 3954
rect 858 3888 868 3954
rect 342 3878 868 3888
rect 970 3858 1500 3868
rect 970 3792 980 3858
rect 1490 3792 1500 3858
rect 970 3782 1500 3792
rect 342 3762 868 3772
rect 342 3696 352 3762
rect 858 3696 868 3762
rect 342 3686 868 3696
rect 970 3666 1500 3676
rect 970 3600 980 3666
rect 1490 3600 1500 3666
rect 970 3590 1500 3600
rect 342 3570 868 3580
rect 342 3504 352 3570
rect 858 3504 868 3570
rect 342 3494 868 3504
rect 970 3474 1500 3484
rect 970 3408 980 3474
rect 1490 3408 1500 3474
rect 970 3398 1500 3408
rect 342 3378 868 3388
rect 342 3312 352 3378
rect 858 3312 868 3378
rect 342 3302 868 3312
rect 970 3282 1500 3292
rect 970 3216 980 3282
rect 1490 3216 1500 3282
rect 970 3206 1500 3216
rect 342 3186 868 3196
rect 342 3120 352 3186
rect 858 3120 868 3186
rect 342 3110 868 3120
rect 970 3090 1500 3100
rect 970 3024 980 3090
rect 1490 3024 1500 3090
rect 970 3014 1500 3024
rect 342 2994 868 3004
rect 342 2928 352 2994
rect 858 2928 868 2994
rect 342 2918 868 2928
rect 970 2898 1500 2908
rect 970 2832 980 2898
rect 1490 2832 1500 2898
rect 970 2822 1500 2832
rect 342 2802 868 2812
rect 342 2736 352 2802
rect 858 2736 868 2802
rect 342 2726 868 2736
rect 970 2706 1500 2716
rect 970 2640 980 2706
rect 1490 2640 1500 2706
rect 970 2630 1500 2640
rect 342 2610 868 2620
rect 342 2544 352 2610
rect 858 2544 868 2610
rect 342 2534 868 2544
rect 970 2514 1500 2524
rect 970 2448 980 2514
rect 1490 2448 1500 2514
rect 970 2438 1500 2448
rect 342 2418 868 2428
rect 342 2352 352 2418
rect 858 2352 868 2418
rect 342 2342 868 2352
rect 970 2322 1500 2332
rect 970 2256 980 2322
rect 1490 2256 1500 2322
rect 970 2246 1500 2256
rect 342 2226 868 2236
rect 342 2160 352 2226
rect 858 2160 868 2226
rect 342 2150 868 2160
rect 970 2130 1500 2140
rect 970 2064 980 2130
rect 1490 2064 1500 2130
rect 970 2054 1500 2064
rect 342 2034 868 2044
rect 342 1968 352 2034
rect 858 1968 868 2034
rect 342 1958 868 1968
rect 970 1938 1500 1948
rect 970 1872 980 1938
rect 1490 1872 1500 1938
rect 970 1862 1500 1872
rect 342 1842 868 1852
rect 342 1776 352 1842
rect 858 1776 868 1842
rect 342 1766 868 1776
rect 970 1746 1500 1756
rect 970 1680 980 1746
rect 1490 1680 1500 1746
rect 970 1670 1500 1680
rect 342 1650 868 1660
rect 342 1584 352 1650
rect 858 1584 868 1650
rect 342 1574 868 1584
rect 970 1554 1500 1564
rect 970 1488 980 1554
rect 1490 1488 1500 1554
rect 970 1478 1500 1488
rect 342 1458 868 1468
rect 342 1392 352 1458
rect 858 1392 868 1458
rect 342 1382 868 1392
rect 970 1362 1500 1372
rect 970 1296 980 1362
rect 1490 1296 1500 1362
rect 970 1286 1500 1296
rect 342 1266 868 1276
rect 342 1200 352 1266
rect 858 1200 868 1266
rect 342 1190 868 1200
rect 970 1170 1500 1180
rect 970 1104 980 1170
rect 1490 1104 1500 1170
rect 970 1094 1500 1104
rect 342 1074 868 1084
rect 342 1008 352 1074
rect 858 1008 868 1074
rect 342 998 868 1008
rect 970 978 1500 988
rect 970 912 980 978
rect 1490 912 1500 978
rect 970 902 1500 912
rect 342 882 868 892
rect 342 816 352 882
rect 858 816 868 882
rect 342 806 868 816
rect 970 786 1500 796
rect 970 720 980 786
rect 1490 720 1500 786
rect 970 710 1500 720
rect 342 690 868 700
rect 342 624 352 690
rect 858 624 868 690
rect 342 614 868 624
<< via3 >>
rect 132 22222 1706 22286
rect 352 21868 858 21934
rect 352 21744 858 21810
rect 980 21648 1490 21714
rect 352 21552 858 21618
rect 980 21456 1490 21522
rect 352 21360 858 21426
rect 980 21264 1490 21330
rect 352 21168 858 21234
rect 980 21072 1490 21138
rect 352 20976 858 21042
rect 980 20880 1490 20946
rect 352 20784 858 20850
rect 980 20688 1490 20754
rect 352 20592 858 20658
rect 980 20496 1490 20562
rect 352 20400 858 20466
rect 980 20304 1490 20370
rect 352 20208 858 20274
rect 980 20112 1490 20178
rect 352 20016 858 20082
rect 980 19920 1490 19986
rect 352 19824 858 19890
rect 980 19728 1490 19794
rect 352 19632 858 19698
rect 980 19536 1490 19602
rect 352 19440 858 19506
rect 980 19344 1490 19410
rect 352 19248 858 19314
rect 980 19152 1490 19218
rect 352 19056 858 19122
rect 980 18960 1490 19026
rect 352 18864 858 18930
rect 980 18768 1490 18834
rect 352 18672 858 18738
rect 980 18576 1490 18642
rect 352 18480 858 18546
rect 980 18384 1490 18450
rect 352 18288 858 18354
rect 980 18192 1490 18258
rect 352 18096 858 18162
rect 980 18000 1490 18066
rect 352 17904 858 17970
rect 980 17808 1490 17874
rect 352 17712 858 17778
rect 980 17616 1490 17682
rect 352 17520 858 17586
rect 980 17424 1490 17490
rect 352 17328 858 17394
rect 980 17232 1490 17298
rect 352 17136 858 17202
rect 980 17040 1490 17106
rect 352 16944 858 17010
rect 980 16848 1490 16914
rect 352 16752 858 16818
rect 980 16656 1490 16722
rect 352 16560 858 16626
rect 980 16464 1490 16530
rect 352 16368 858 16434
rect 980 16272 1490 16338
rect 352 16176 858 16242
rect 980 16080 1490 16146
rect 352 15984 858 16050
rect 980 15888 1490 15954
rect 352 15792 858 15858
rect 980 15696 1490 15762
rect 352 15600 858 15666
rect 980 15504 1490 15570
rect 352 15408 858 15474
rect 980 15312 1490 15378
rect 352 15216 858 15282
rect 980 15120 1490 15186
rect 352 15024 858 15090
rect 980 14928 1490 14994
rect 352 14832 858 14898
rect 980 14736 1490 14802
rect 352 14640 858 14706
rect 980 14544 1490 14610
rect 352 14448 858 14514
rect 980 14352 1490 14418
rect 352 14256 858 14322
rect 980 14160 1490 14226
rect 352 14064 858 14130
rect 980 13968 1490 14034
rect 352 13872 858 13938
rect 980 13776 1490 13842
rect 352 13680 858 13746
rect 980 13584 1490 13650
rect 352 13488 858 13554
rect 980 13392 1490 13458
rect 352 13296 858 13362
rect 980 13200 1490 13266
rect 352 13104 858 13170
rect 980 13008 1490 13074
rect 352 12912 858 12978
rect 980 12816 1490 12882
rect 352 12720 858 12786
rect 980 12624 1490 12690
rect 352 12528 858 12594
rect 980 12432 1490 12498
rect 352 12336 858 12402
rect 980 12240 1490 12306
rect 352 12144 858 12210
rect 980 12048 1490 12114
rect 352 11952 858 12018
rect 980 11856 1490 11922
rect 352 11760 858 11826
rect 980 11664 1490 11730
rect 352 11568 858 11634
rect 980 11472 1490 11538
rect 352 11376 858 11442
rect 980 11280 1490 11346
rect 352 11184 858 11250
rect 980 11088 1490 11154
rect 352 10992 858 11058
rect 980 10896 1490 10962
rect 352 10800 858 10866
rect 980 10704 1490 10770
rect 352 10608 858 10674
rect 980 10512 1490 10578
rect 352 10416 858 10482
rect 980 10320 1490 10386
rect 352 10224 858 10290
rect 980 10128 1490 10194
rect 352 10032 858 10098
rect 980 9936 1490 10002
rect 352 9840 858 9906
rect 980 9744 1490 9810
rect 352 9648 858 9714
rect 980 9552 1490 9618
rect 352 9456 858 9522
rect 980 9360 1490 9426
rect 352 9264 858 9330
rect 980 9168 1490 9234
rect 352 9072 858 9138
rect 980 8976 1490 9042
rect 352 8880 858 8946
rect 980 8784 1490 8850
rect 352 8688 858 8754
rect 980 8592 1490 8658
rect 352 8496 858 8562
rect 980 8400 1490 8466
rect 352 8304 858 8370
rect 980 8208 1490 8274
rect 352 8112 858 8178
rect 980 8016 1490 8082
rect 352 7920 858 7986
rect 980 7824 1490 7890
rect 352 7728 858 7794
rect 980 7632 1490 7698
rect 352 7536 858 7602
rect 980 7440 1490 7506
rect 352 7344 858 7410
rect 980 7248 1490 7314
rect 352 7152 858 7218
rect 980 7056 1490 7122
rect 352 6960 858 7026
rect 980 6864 1490 6930
rect 352 6768 858 6834
rect 980 6672 1490 6738
rect 352 6576 858 6642
rect 980 6480 1490 6546
rect 352 6384 858 6450
rect 980 6288 1490 6354
rect 352 6192 858 6258
rect 980 6096 1490 6162
rect 352 6000 858 6066
rect 980 5904 1490 5970
rect 352 5808 858 5874
rect 980 5712 1490 5778
rect 352 5616 858 5682
rect 980 5520 1490 5586
rect 352 5424 858 5490
rect 980 5328 1490 5394
rect 352 5232 858 5298
rect 980 5136 1490 5202
rect 352 5040 858 5106
rect 980 4944 1490 5010
rect 352 4848 858 4914
rect 980 4752 1490 4818
rect 352 4656 858 4722
rect 980 4560 1490 4626
rect 352 4464 858 4530
rect 980 4368 1490 4434
rect 352 4272 858 4338
rect 980 4176 1490 4242
rect 352 4080 858 4146
rect 980 3984 1490 4050
rect 352 3888 858 3954
rect 980 3792 1490 3858
rect 352 3696 858 3762
rect 980 3600 1490 3666
rect 352 3504 858 3570
rect 980 3408 1490 3474
rect 352 3312 858 3378
rect 980 3216 1490 3282
rect 352 3120 858 3186
rect 980 3024 1490 3090
rect 352 2928 858 2994
rect 980 2832 1490 2898
rect 352 2736 858 2802
rect 980 2640 1490 2706
rect 352 2544 858 2610
rect 980 2448 1490 2514
rect 352 2352 858 2418
rect 980 2256 1490 2322
rect 352 2160 858 2226
rect 980 2064 1490 2130
rect 352 1968 858 2034
rect 980 1872 1490 1938
rect 352 1776 858 1842
rect 980 1680 1490 1746
rect 352 1584 858 1650
rect 980 1488 1490 1554
rect 352 1392 858 1458
rect 980 1296 1490 1362
rect 352 1200 858 1266
rect 980 1104 1490 1170
rect 352 1008 858 1074
rect 980 912 1490 978
rect 352 816 858 882
rect 980 720 1490 786
rect 352 624 858 690
<< metal4 >>
rect 0 22286 1840 22304
rect 0 22222 132 22286
rect 1706 22222 1840 22286
rect 0 22204 1840 22222
rect 0 0 240 22000
rect 340 21934 870 22000
rect 340 21868 352 21934
rect 858 21868 870 21934
rect 340 21810 870 21868
rect 340 21744 352 21810
rect 858 21744 870 21810
rect 340 21618 870 21744
rect 340 21552 352 21618
rect 858 21552 870 21618
rect 340 21426 870 21552
rect 340 21360 352 21426
rect 858 21360 870 21426
rect 340 21234 870 21360
rect 340 21168 352 21234
rect 858 21168 870 21234
rect 340 21042 870 21168
rect 340 20976 352 21042
rect 858 20976 870 21042
rect 340 20850 870 20976
rect 340 20784 352 20850
rect 858 20784 870 20850
rect 340 20658 870 20784
rect 340 20592 352 20658
rect 858 20592 870 20658
rect 340 20466 870 20592
rect 340 20400 352 20466
rect 858 20400 870 20466
rect 340 20274 870 20400
rect 340 20208 352 20274
rect 858 20208 870 20274
rect 340 20082 870 20208
rect 340 20016 352 20082
rect 858 20016 870 20082
rect 340 19890 870 20016
rect 340 19824 352 19890
rect 858 19824 870 19890
rect 340 19698 870 19824
rect 340 19632 352 19698
rect 858 19632 870 19698
rect 340 19506 870 19632
rect 340 19440 352 19506
rect 858 19440 870 19506
rect 340 19314 870 19440
rect 340 19248 352 19314
rect 858 19248 870 19314
rect 340 19122 870 19248
rect 340 19056 352 19122
rect 858 19056 870 19122
rect 340 18930 870 19056
rect 340 18864 352 18930
rect 858 18864 870 18930
rect 340 18738 870 18864
rect 340 18672 352 18738
rect 858 18672 870 18738
rect 340 18546 870 18672
rect 340 18480 352 18546
rect 858 18480 870 18546
rect 340 18354 870 18480
rect 340 18288 352 18354
rect 858 18288 870 18354
rect 340 18162 870 18288
rect 340 18096 352 18162
rect 858 18096 870 18162
rect 340 17970 870 18096
rect 340 17904 352 17970
rect 858 17904 870 17970
rect 340 17778 870 17904
rect 340 17712 352 17778
rect 858 17712 870 17778
rect 340 17586 870 17712
rect 340 17520 352 17586
rect 858 17520 870 17586
rect 340 17394 870 17520
rect 340 17328 352 17394
rect 858 17328 870 17394
rect 340 17202 870 17328
rect 340 17136 352 17202
rect 858 17136 870 17202
rect 340 17010 870 17136
rect 340 16944 352 17010
rect 858 16944 870 17010
rect 340 16818 870 16944
rect 340 16752 352 16818
rect 858 16752 870 16818
rect 340 16626 870 16752
rect 340 16560 352 16626
rect 858 16560 870 16626
rect 340 16434 870 16560
rect 340 16368 352 16434
rect 858 16368 870 16434
rect 340 16242 870 16368
rect 340 16176 352 16242
rect 858 16176 870 16242
rect 340 16050 870 16176
rect 340 15984 352 16050
rect 858 15984 870 16050
rect 340 15858 870 15984
rect 340 15792 352 15858
rect 858 15792 870 15858
rect 340 15666 870 15792
rect 340 15600 352 15666
rect 858 15600 870 15666
rect 340 15474 870 15600
rect 340 15408 352 15474
rect 858 15408 870 15474
rect 340 15282 870 15408
rect 340 15216 352 15282
rect 858 15216 870 15282
rect 340 15090 870 15216
rect 340 15024 352 15090
rect 858 15024 870 15090
rect 340 14898 870 15024
rect 340 14832 352 14898
rect 858 14832 870 14898
rect 340 14706 870 14832
rect 340 14640 352 14706
rect 858 14640 870 14706
rect 340 14514 870 14640
rect 340 14448 352 14514
rect 858 14448 870 14514
rect 340 14322 870 14448
rect 340 14256 352 14322
rect 858 14256 870 14322
rect 340 14130 870 14256
rect 340 14064 352 14130
rect 858 14064 870 14130
rect 340 13938 870 14064
rect 340 13872 352 13938
rect 858 13872 870 13938
rect 340 13746 870 13872
rect 340 13680 352 13746
rect 858 13680 870 13746
rect 340 13554 870 13680
rect 340 13488 352 13554
rect 858 13488 870 13554
rect 340 13362 870 13488
rect 340 13296 352 13362
rect 858 13296 870 13362
rect 340 13170 870 13296
rect 340 13104 352 13170
rect 858 13104 870 13170
rect 340 12978 870 13104
rect 340 12912 352 12978
rect 858 12912 870 12978
rect 340 12786 870 12912
rect 340 12720 352 12786
rect 858 12720 870 12786
rect 340 12594 870 12720
rect 340 12528 352 12594
rect 858 12528 870 12594
rect 340 12402 870 12528
rect 340 12336 352 12402
rect 858 12336 870 12402
rect 340 12210 870 12336
rect 340 12144 352 12210
rect 858 12144 870 12210
rect 340 12018 870 12144
rect 340 11952 352 12018
rect 858 11952 870 12018
rect 340 11826 870 11952
rect 340 11760 352 11826
rect 858 11760 870 11826
rect 340 11634 870 11760
rect 340 11568 352 11634
rect 858 11568 870 11634
rect 340 11442 870 11568
rect 340 11376 352 11442
rect 858 11376 870 11442
rect 340 11250 870 11376
rect 340 11184 352 11250
rect 858 11184 870 11250
rect 340 11058 870 11184
rect 340 10992 352 11058
rect 858 10992 870 11058
rect 340 10866 870 10992
rect 340 10800 352 10866
rect 858 10800 870 10866
rect 340 10674 870 10800
rect 340 10608 352 10674
rect 858 10608 870 10674
rect 340 10482 870 10608
rect 340 10416 352 10482
rect 858 10416 870 10482
rect 340 10290 870 10416
rect 340 10224 352 10290
rect 858 10224 870 10290
rect 340 10098 870 10224
rect 340 10032 352 10098
rect 858 10032 870 10098
rect 340 9906 870 10032
rect 340 9840 352 9906
rect 858 9840 870 9906
rect 340 9714 870 9840
rect 340 9648 352 9714
rect 858 9648 870 9714
rect 340 9522 870 9648
rect 340 9456 352 9522
rect 858 9456 870 9522
rect 340 9330 870 9456
rect 340 9264 352 9330
rect 858 9264 870 9330
rect 340 9138 870 9264
rect 340 9072 352 9138
rect 858 9072 870 9138
rect 340 8946 870 9072
rect 340 8880 352 8946
rect 858 8880 870 8946
rect 340 8754 870 8880
rect 340 8688 352 8754
rect 858 8688 870 8754
rect 340 8562 870 8688
rect 340 8496 352 8562
rect 858 8496 870 8562
rect 340 8370 870 8496
rect 340 8304 352 8370
rect 858 8304 870 8370
rect 340 8178 870 8304
rect 340 8112 352 8178
rect 858 8112 870 8178
rect 340 7986 870 8112
rect 340 7920 352 7986
rect 858 7920 870 7986
rect 340 7794 870 7920
rect 340 7728 352 7794
rect 858 7728 870 7794
rect 340 7602 870 7728
rect 340 7536 352 7602
rect 858 7536 870 7602
rect 340 7410 870 7536
rect 340 7344 352 7410
rect 858 7344 870 7410
rect 340 7218 870 7344
rect 340 7152 352 7218
rect 858 7152 870 7218
rect 340 7026 870 7152
rect 340 6960 352 7026
rect 858 6960 870 7026
rect 340 6834 870 6960
rect 340 6768 352 6834
rect 858 6768 870 6834
rect 340 6642 870 6768
rect 340 6576 352 6642
rect 858 6576 870 6642
rect 340 6450 870 6576
rect 340 6384 352 6450
rect 858 6384 870 6450
rect 340 6258 870 6384
rect 340 6192 352 6258
rect 858 6192 870 6258
rect 340 6066 870 6192
rect 340 6000 352 6066
rect 858 6000 870 6066
rect 340 5874 870 6000
rect 340 5808 352 5874
rect 858 5808 870 5874
rect 340 5682 870 5808
rect 340 5616 352 5682
rect 858 5616 870 5682
rect 340 5490 870 5616
rect 340 5424 352 5490
rect 858 5424 870 5490
rect 340 5298 870 5424
rect 340 5232 352 5298
rect 858 5232 870 5298
rect 340 5106 870 5232
rect 340 5040 352 5106
rect 858 5040 870 5106
rect 340 4914 870 5040
rect 340 4848 352 4914
rect 858 4848 870 4914
rect 340 4722 870 4848
rect 340 4656 352 4722
rect 858 4656 870 4722
rect 340 4530 870 4656
rect 340 4464 352 4530
rect 858 4464 870 4530
rect 340 4338 870 4464
rect 340 4272 352 4338
rect 858 4272 870 4338
rect 340 4146 870 4272
rect 340 4080 352 4146
rect 858 4080 870 4146
rect 340 3954 870 4080
rect 340 3888 352 3954
rect 858 3888 870 3954
rect 340 3762 870 3888
rect 340 3696 352 3762
rect 858 3696 870 3762
rect 340 3570 870 3696
rect 340 3504 352 3570
rect 858 3504 870 3570
rect 340 3378 870 3504
rect 340 3312 352 3378
rect 858 3312 870 3378
rect 340 3186 870 3312
rect 340 3120 352 3186
rect 858 3120 870 3186
rect 340 2994 870 3120
rect 340 2928 352 2994
rect 858 2928 870 2994
rect 340 2802 870 2928
rect 340 2736 352 2802
rect 858 2736 870 2802
rect 340 2610 870 2736
rect 340 2544 352 2610
rect 858 2544 870 2610
rect 340 2418 870 2544
rect 340 2352 352 2418
rect 858 2352 870 2418
rect 340 2226 870 2352
rect 340 2160 352 2226
rect 858 2160 870 2226
rect 340 2089 870 2160
rect 970 21714 1500 22000
rect 970 21648 980 21714
rect 1490 21648 1500 21714
rect 970 21522 1500 21648
rect 970 21456 980 21522
rect 1490 21456 1500 21522
rect 970 21330 1500 21456
rect 970 21264 980 21330
rect 1490 21264 1500 21330
rect 970 21138 1500 21264
rect 970 21072 980 21138
rect 1490 21072 1500 21138
rect 970 20946 1500 21072
rect 970 20880 980 20946
rect 1490 20880 1500 20946
rect 970 20754 1500 20880
rect 970 20688 980 20754
rect 1490 20688 1500 20754
rect 970 20562 1500 20688
rect 970 20496 980 20562
rect 1490 20496 1500 20562
rect 970 20370 1500 20496
rect 970 20304 980 20370
rect 1490 20304 1500 20370
rect 970 20178 1500 20304
rect 970 20112 980 20178
rect 1490 20112 1500 20178
rect 970 19986 1500 20112
rect 970 19920 980 19986
rect 1490 19920 1500 19986
rect 970 19794 1500 19920
rect 970 19728 980 19794
rect 1490 19728 1500 19794
rect 970 19602 1500 19728
rect 970 19536 980 19602
rect 1490 19536 1500 19602
rect 970 19410 1500 19536
rect 970 19344 980 19410
rect 1490 19344 1500 19410
rect 970 19218 1500 19344
rect 970 19152 980 19218
rect 1490 19152 1500 19218
rect 970 19026 1500 19152
rect 970 18960 980 19026
rect 1490 18960 1500 19026
rect 970 18834 1500 18960
rect 970 18768 980 18834
rect 1490 18768 1500 18834
rect 970 18642 1500 18768
rect 970 18576 980 18642
rect 1490 18576 1500 18642
rect 970 18450 1500 18576
rect 970 18384 980 18450
rect 1490 18384 1500 18450
rect 970 18258 1500 18384
rect 970 18192 980 18258
rect 1490 18192 1500 18258
rect 970 18066 1500 18192
rect 970 18000 980 18066
rect 1490 18000 1500 18066
rect 970 17874 1500 18000
rect 970 17808 980 17874
rect 1490 17808 1500 17874
rect 970 17682 1500 17808
rect 970 17616 980 17682
rect 1490 17616 1500 17682
rect 970 17490 1500 17616
rect 970 17424 980 17490
rect 1490 17424 1500 17490
rect 970 17298 1500 17424
rect 970 17232 980 17298
rect 1490 17232 1500 17298
rect 970 17106 1500 17232
rect 970 17040 980 17106
rect 1490 17040 1500 17106
rect 970 16914 1500 17040
rect 970 16848 980 16914
rect 1490 16848 1500 16914
rect 970 16722 1500 16848
rect 970 16656 980 16722
rect 1490 16656 1500 16722
rect 970 16530 1500 16656
rect 970 16464 980 16530
rect 1490 16464 1500 16530
rect 970 16338 1500 16464
rect 970 16272 980 16338
rect 1490 16272 1500 16338
rect 970 16146 1500 16272
rect 970 16080 980 16146
rect 1490 16080 1500 16146
rect 970 15954 1500 16080
rect 970 15888 980 15954
rect 1490 15888 1500 15954
rect 970 15762 1500 15888
rect 970 15696 980 15762
rect 1490 15696 1500 15762
rect 970 15570 1500 15696
rect 970 15504 980 15570
rect 1490 15504 1500 15570
rect 970 15378 1500 15504
rect 970 15312 980 15378
rect 1490 15312 1500 15378
rect 970 15186 1500 15312
rect 970 15120 980 15186
rect 1490 15120 1500 15186
rect 970 14994 1500 15120
rect 970 14928 980 14994
rect 1490 14928 1500 14994
rect 970 14802 1500 14928
rect 970 14736 980 14802
rect 1490 14736 1500 14802
rect 970 14610 1500 14736
rect 970 14544 980 14610
rect 1490 14544 1500 14610
rect 970 14418 1500 14544
rect 970 14352 980 14418
rect 1490 14352 1500 14418
rect 970 14226 1500 14352
rect 970 14160 980 14226
rect 1490 14160 1500 14226
rect 970 14034 1500 14160
rect 970 13968 980 14034
rect 1490 13968 1500 14034
rect 970 13842 1500 13968
rect 970 13776 980 13842
rect 1490 13776 1500 13842
rect 970 13650 1500 13776
rect 970 13584 980 13650
rect 1490 13584 1500 13650
rect 970 13458 1500 13584
rect 970 13392 980 13458
rect 1490 13392 1500 13458
rect 970 13266 1500 13392
rect 970 13200 980 13266
rect 1490 13200 1500 13266
rect 970 13074 1500 13200
rect 970 13008 980 13074
rect 1490 13008 1500 13074
rect 970 12882 1500 13008
rect 970 12816 980 12882
rect 1490 12816 1500 12882
rect 970 12690 1500 12816
rect 970 12624 980 12690
rect 1490 12624 1500 12690
rect 970 12498 1500 12624
rect 970 12432 980 12498
rect 1490 12432 1500 12498
rect 970 12306 1500 12432
rect 970 12240 980 12306
rect 1490 12240 1500 12306
rect 970 12114 1500 12240
rect 970 12048 980 12114
rect 1490 12048 1500 12114
rect 970 11922 1500 12048
rect 970 11856 980 11922
rect 1490 11856 1500 11922
rect 970 11730 1500 11856
rect 970 11664 980 11730
rect 1490 11664 1500 11730
rect 970 11538 1500 11664
rect 970 11472 980 11538
rect 1490 11472 1500 11538
rect 970 11346 1500 11472
rect 970 11280 980 11346
rect 1490 11280 1500 11346
rect 970 11154 1500 11280
rect 970 11088 980 11154
rect 1490 11088 1500 11154
rect 970 10962 1500 11088
rect 970 10896 980 10962
rect 1490 10896 1500 10962
rect 970 10770 1500 10896
rect 970 10704 980 10770
rect 1490 10704 1500 10770
rect 970 10578 1500 10704
rect 970 10512 980 10578
rect 1490 10512 1500 10578
rect 970 10386 1500 10512
rect 970 10320 980 10386
rect 1490 10320 1500 10386
rect 970 10194 1500 10320
rect 970 10128 980 10194
rect 1490 10128 1500 10194
rect 970 10002 1500 10128
rect 970 9936 980 10002
rect 1490 9936 1500 10002
rect 970 9810 1500 9936
rect 970 9744 980 9810
rect 1490 9744 1500 9810
rect 970 9618 1500 9744
rect 970 9552 980 9618
rect 1490 9552 1500 9618
rect 970 9426 1500 9552
rect 970 9360 980 9426
rect 1490 9360 1500 9426
rect 970 9234 1500 9360
rect 970 9168 980 9234
rect 1490 9168 1500 9234
rect 970 9042 1500 9168
rect 970 8976 980 9042
rect 1490 8976 1500 9042
rect 970 8850 1500 8976
rect 970 8784 980 8850
rect 1490 8784 1500 8850
rect 970 8658 1500 8784
rect 970 8592 980 8658
rect 1490 8592 1500 8658
rect 970 8466 1500 8592
rect 970 8400 980 8466
rect 1490 8400 1500 8466
rect 970 8274 1500 8400
rect 970 8208 980 8274
rect 1490 8208 1500 8274
rect 970 8082 1500 8208
rect 970 8016 980 8082
rect 1490 8016 1500 8082
rect 970 7890 1500 8016
rect 970 7824 980 7890
rect 1490 7824 1500 7890
rect 970 7698 1500 7824
rect 970 7632 980 7698
rect 1490 7632 1500 7698
rect 970 7506 1500 7632
rect 970 7440 980 7506
rect 1490 7440 1500 7506
rect 970 7314 1500 7440
rect 970 7248 980 7314
rect 1490 7248 1500 7314
rect 970 7122 1500 7248
rect 970 7056 980 7122
rect 1490 7056 1500 7122
rect 970 6930 1500 7056
rect 970 6864 980 6930
rect 1490 6864 1500 6930
rect 970 6738 1500 6864
rect 970 6672 980 6738
rect 1490 6672 1500 6738
rect 970 6546 1500 6672
rect 970 6480 980 6546
rect 1490 6480 1500 6546
rect 970 6354 1500 6480
rect 970 6288 980 6354
rect 1490 6288 1500 6354
rect 970 6162 1500 6288
rect 970 6096 980 6162
rect 1490 6096 1500 6162
rect 970 5970 1500 6096
rect 970 5904 980 5970
rect 1490 5904 1500 5970
rect 970 5778 1500 5904
rect 970 5712 980 5778
rect 1490 5712 1500 5778
rect 970 5586 1500 5712
rect 970 5520 980 5586
rect 1490 5520 1500 5586
rect 970 5394 1500 5520
rect 970 5328 980 5394
rect 1490 5328 1500 5394
rect 970 5202 1500 5328
rect 970 5136 980 5202
rect 1490 5136 1500 5202
rect 970 5010 1500 5136
rect 970 4944 980 5010
rect 1490 4944 1500 5010
rect 970 4818 1500 4944
rect 970 4752 980 4818
rect 1490 4752 1500 4818
rect 970 4626 1500 4752
rect 970 4560 980 4626
rect 1490 4560 1500 4626
rect 970 4434 1500 4560
rect 970 4368 980 4434
rect 1490 4368 1500 4434
rect 970 4242 1500 4368
rect 970 4176 980 4242
rect 1490 4176 1500 4242
rect 970 4050 1500 4176
rect 970 3984 980 4050
rect 1490 3984 1500 4050
rect 970 3858 1500 3984
rect 970 3792 980 3858
rect 1490 3792 1500 3858
rect 970 3666 1500 3792
rect 970 3600 980 3666
rect 1490 3600 1500 3666
rect 970 3474 1500 3600
rect 970 3408 980 3474
rect 1490 3408 1500 3474
rect 970 3282 1500 3408
rect 970 3216 980 3282
rect 1490 3216 1500 3282
rect 970 3090 1500 3216
rect 970 3024 980 3090
rect 1490 3024 1500 3090
rect 970 2898 1500 3024
rect 970 2832 980 2898
rect 1490 2832 1500 2898
rect 970 2706 1500 2832
rect 970 2640 980 2706
rect 1490 2640 1500 2706
rect 970 2514 1500 2640
rect 970 2448 980 2514
rect 1490 2448 1500 2514
rect 970 2322 1500 2448
rect 970 2256 980 2322
rect 1490 2256 1500 2322
rect 970 2130 1500 2256
rect 339 2034 871 2089
rect 339 2023 352 2034
rect 340 1968 352 2023
rect 858 2023 871 2034
rect 970 2064 980 2130
rect 1490 2064 1500 2130
rect 858 1968 870 2023
rect 340 1899 870 1968
rect 970 1938 1500 2064
rect 339 1842 871 1899
rect 339 1833 352 1842
rect 340 1776 352 1833
rect 858 1833 871 1842
rect 970 1872 980 1938
rect 1490 1872 1500 1938
rect 858 1776 870 1833
rect 340 1705 870 1776
rect 970 1746 1500 1872
rect 339 1650 871 1705
rect 339 1639 352 1650
rect 340 1584 352 1639
rect 858 1639 871 1650
rect 970 1680 980 1746
rect 1490 1680 1500 1746
rect 858 1584 870 1639
rect 340 1515 870 1584
rect 970 1554 1500 1680
rect 339 1458 871 1515
rect 339 1449 352 1458
rect 340 1392 352 1449
rect 858 1449 871 1458
rect 970 1488 980 1554
rect 1490 1488 1500 1554
rect 858 1392 870 1449
rect 340 1323 870 1392
rect 970 1362 1500 1488
rect 339 1266 871 1323
rect 339 1257 352 1266
rect 340 1200 352 1257
rect 858 1257 871 1266
rect 970 1296 980 1362
rect 1490 1296 1500 1362
rect 858 1200 870 1257
rect 340 1129 870 1200
rect 970 1170 1500 1296
rect 339 1074 871 1129
rect 339 1063 352 1074
rect 340 1008 352 1063
rect 858 1063 871 1074
rect 970 1104 980 1170
rect 1490 1104 1500 1170
rect 858 1008 870 1063
rect 340 939 870 1008
rect 970 978 1500 1104
rect 339 882 871 939
rect 339 873 352 882
rect 340 816 352 873
rect 858 873 871 882
rect 970 912 980 978
rect 1490 912 1500 978
rect 858 816 870 873
rect 340 747 870 816
rect 970 786 1500 912
rect 339 690 871 747
rect 339 681 352 690
rect 340 624 352 681
rect 858 681 871 690
rect 970 720 980 786
rect 1490 720 1500 786
rect 858 624 870 681
rect 340 0 870 624
rect 970 0 1500 720
rect 1600 0 1840 22000
<< labels >>
rlabel metal4 0 0 240 22000 1 VGND
port 1 n ground input
rlabel metal4 1600 0 1840 22000 1 VGND
port 1 n ground input
rlabel metal4 340 0 870 22000 1 VPWR
port 2 n power input
rlabel metal4 970 0 1500 22000 1 GPWR
port 3 n power output
rlabel metal4 0 22204 1840 22304 1 ctrl
port 4 n signal input
<< properties >>
string FIXED_BBOX 0 0 1840 22304
<< end >>
