magic
tech sky130A
magscale 1 2
timestamp 1718383489
<< metal3 >>
rect 340 3994 2660 4000
rect 340 6 341 3994
rect 579 6 2660 3994
rect 340 0 2660 6
<< via3 >>
rect 341 6 579 3994
<< mimcap >>
rect 640 3880 2600 3940
rect 640 120 740 3880
rect 1610 120 2600 3880
rect 640 60 2600 120
<< mimcapcontact >>
rect 740 120 1610 3880
<< metal4 >>
rect 0 0 240 4000
rect 340 3994 580 4000
rect 340 6 341 3994
rect 579 6 580 3994
rect 340 0 580 6
rect 680 3880 1670 4000
rect 680 120 740 3880
rect 1610 120 1670 3880
rect 680 0 1670 120
rect 1770 0 2760 4000
<< end >>
