module vssd1_connection ();
endmodule