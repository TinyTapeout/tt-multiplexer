magic
tech sky130A
magscale 1 2
timestamp 1718204978
<< nwell >>
rect 0 0 1780 43994
<< pmos >>
rect 130 43783 1580 43813
rect 130 43697 1580 43727
rect 130 43611 1580 43641
rect 130 43525 1580 43555
rect 130 43439 1580 43469
rect 130 43353 1580 43383
rect 130 43267 1580 43297
rect 130 43181 1580 43211
rect 130 43095 1580 43125
rect 130 43009 1580 43039
rect 130 42923 1580 42953
rect 130 42837 1580 42867
rect 130 42751 1580 42781
rect 130 42665 1580 42695
rect 130 42579 1580 42609
rect 130 42493 1580 42523
rect 130 42407 1580 42437
rect 130 42321 1580 42351
rect 130 42235 1580 42265
rect 130 42149 1580 42179
rect 130 42063 1580 42093
rect 130 41977 1580 42007
rect 130 41891 1580 41921
rect 130 41805 1580 41835
rect 130 41719 1580 41749
rect 130 41633 1580 41663
rect 130 41547 1580 41577
rect 130 41461 1580 41491
rect 130 41375 1580 41405
rect 130 41289 1580 41319
rect 130 41203 1580 41233
rect 130 41117 1580 41147
rect 130 41031 1580 41061
rect 130 40945 1580 40975
rect 130 40859 1580 40889
rect 130 40773 1580 40803
rect 130 40687 1580 40717
rect 130 40601 1580 40631
rect 130 40515 1580 40545
rect 130 40429 1580 40459
rect 130 40343 1580 40373
rect 130 40257 1580 40287
rect 130 40171 1580 40201
rect 130 40085 1580 40115
rect 130 39999 1580 40029
rect 130 39913 1580 39943
rect 130 39827 1580 39857
rect 130 39741 1580 39771
rect 130 39655 1580 39685
rect 130 39569 1580 39599
rect 130 39483 1580 39513
rect 130 39397 1580 39427
rect 130 39311 1580 39341
rect 130 39225 1580 39255
rect 130 39139 1580 39169
rect 130 39053 1580 39083
rect 130 38967 1580 38997
rect 130 38881 1580 38911
rect 130 38795 1580 38825
rect 130 38709 1580 38739
rect 130 38623 1580 38653
rect 130 38537 1580 38567
rect 130 38451 1580 38481
rect 130 38365 1580 38395
rect 130 38279 1580 38309
rect 130 38193 1580 38223
rect 130 38107 1580 38137
rect 130 38021 1580 38051
rect 130 37935 1580 37965
rect 130 37849 1580 37879
rect 130 37763 1580 37793
rect 130 37677 1580 37707
rect 130 37591 1580 37621
rect 130 37505 1580 37535
rect 130 37419 1580 37449
rect 130 37333 1580 37363
rect 130 37247 1580 37277
rect 130 37161 1580 37191
rect 130 37075 1580 37105
rect 130 36989 1580 37019
rect 130 36903 1580 36933
rect 130 36817 1580 36847
rect 130 36731 1580 36761
rect 130 36645 1580 36675
rect 130 36559 1580 36589
rect 130 36473 1580 36503
rect 130 36387 1580 36417
rect 130 36301 1580 36331
rect 130 36215 1580 36245
rect 130 36129 1580 36159
rect 130 36043 1580 36073
rect 130 35957 1580 35987
rect 130 35871 1580 35901
rect 130 35785 1580 35815
rect 130 35699 1580 35729
rect 130 35613 1580 35643
rect 130 35527 1580 35557
rect 130 35441 1580 35471
rect 130 35355 1580 35385
rect 130 35269 1580 35299
rect 130 35183 1580 35213
rect 130 35097 1580 35127
rect 130 35011 1580 35041
rect 130 34925 1580 34955
rect 130 34839 1580 34869
rect 130 34753 1580 34783
rect 130 34667 1580 34697
rect 130 34581 1580 34611
rect 130 34495 1580 34525
rect 130 34409 1580 34439
rect 130 34323 1580 34353
rect 130 34237 1580 34267
rect 130 34151 1580 34181
rect 130 34065 1580 34095
rect 130 33979 1580 34009
rect 130 33893 1580 33923
rect 130 33807 1580 33837
rect 130 33721 1580 33751
rect 130 33635 1580 33665
rect 130 33549 1580 33579
rect 130 33463 1580 33493
rect 130 33377 1580 33407
rect 130 33291 1580 33321
rect 130 33205 1580 33235
rect 130 33119 1580 33149
rect 130 33033 1580 33063
rect 130 32947 1580 32977
rect 130 32861 1580 32891
rect 130 32775 1580 32805
rect 130 32689 1580 32719
rect 130 32603 1580 32633
rect 130 32517 1580 32547
rect 130 32431 1580 32461
rect 130 32345 1580 32375
rect 130 32259 1580 32289
rect 130 32173 1580 32203
rect 130 32087 1580 32117
rect 130 32001 1580 32031
rect 130 31915 1580 31945
rect 130 31829 1580 31859
rect 130 31743 1580 31773
rect 130 31657 1580 31687
rect 130 31571 1580 31601
rect 130 31485 1580 31515
rect 130 31399 1580 31429
rect 130 31313 1580 31343
rect 130 31227 1580 31257
rect 130 31141 1580 31171
rect 130 31055 1580 31085
rect 130 30969 1580 30999
rect 130 30883 1580 30913
rect 130 30797 1580 30827
rect 130 30711 1580 30741
rect 130 30625 1580 30655
rect 130 30539 1580 30569
rect 130 30453 1580 30483
rect 130 30367 1580 30397
rect 130 30281 1580 30311
rect 130 30195 1580 30225
rect 130 30109 1580 30139
rect 130 30023 1580 30053
rect 130 29937 1580 29967
rect 130 29851 1580 29881
rect 130 29765 1580 29795
rect 130 29679 1580 29709
rect 130 29593 1580 29623
rect 130 29507 1580 29537
rect 130 29421 1580 29451
rect 130 29335 1580 29365
rect 130 29249 1580 29279
rect 130 29163 1580 29193
rect 130 29077 1580 29107
rect 130 28991 1580 29021
rect 130 28905 1580 28935
rect 130 28819 1580 28849
rect 130 28733 1580 28763
rect 130 28647 1580 28677
rect 130 28561 1580 28591
rect 130 28475 1580 28505
rect 130 28389 1580 28419
rect 130 28303 1580 28333
rect 130 28217 1580 28247
rect 130 28131 1580 28161
rect 130 28045 1580 28075
rect 130 27959 1580 27989
rect 130 27873 1580 27903
rect 130 27787 1580 27817
rect 130 27701 1580 27731
rect 130 27615 1580 27645
rect 130 27529 1580 27559
rect 130 27443 1580 27473
rect 130 27357 1580 27387
rect 130 27271 1580 27301
rect 130 27185 1580 27215
rect 130 27099 1580 27129
rect 130 27013 1580 27043
rect 130 26927 1580 26957
rect 130 26841 1580 26871
rect 130 26755 1580 26785
rect 130 26669 1580 26699
rect 130 26583 1580 26613
rect 130 26497 1580 26527
rect 130 26411 1580 26441
rect 130 26325 1580 26355
rect 130 26239 1580 26269
rect 130 26153 1580 26183
rect 130 26067 1580 26097
rect 130 25981 1580 26011
rect 130 25895 1580 25925
rect 130 25809 1580 25839
rect 130 25723 1580 25753
rect 130 25637 1580 25667
rect 130 25551 1580 25581
rect 130 25465 1580 25495
rect 130 25379 1580 25409
rect 130 25293 1580 25323
rect 130 25207 1580 25237
rect 130 25121 1580 25151
rect 130 25035 1580 25065
rect 130 24949 1580 24979
rect 130 24863 1580 24893
rect 130 24777 1580 24807
rect 130 24691 1580 24721
rect 130 24605 1580 24635
rect 130 24519 1580 24549
rect 130 24433 1580 24463
rect 130 24347 1580 24377
rect 130 24261 1580 24291
rect 130 24175 1580 24205
rect 130 24089 1580 24119
rect 130 24003 1580 24033
rect 130 23917 1580 23947
rect 130 23831 1580 23861
rect 130 23745 1580 23775
rect 130 23659 1580 23689
rect 130 23573 1580 23603
rect 130 23487 1580 23517
rect 130 23401 1580 23431
rect 130 23315 1580 23345
rect 130 23229 1580 23259
rect 130 23143 1580 23173
rect 130 23057 1580 23087
rect 130 22971 1580 23001
rect 130 22885 1580 22915
rect 130 22799 1580 22829
rect 130 22713 1580 22743
rect 130 22627 1580 22657
rect 130 22541 1580 22571
rect 130 22455 1580 22485
rect 130 22369 1580 22399
rect 130 22283 1580 22313
rect 130 22197 1580 22227
rect 130 22111 1580 22141
rect 130 22025 1580 22055
rect 130 21939 1580 21969
rect 130 21853 1580 21883
rect 130 21767 1580 21797
rect 130 21681 1580 21711
rect 130 21595 1580 21625
rect 130 21509 1580 21539
rect 130 21423 1580 21453
rect 130 21337 1580 21367
rect 130 21251 1580 21281
rect 130 21165 1580 21195
rect 130 21079 1580 21109
rect 130 20993 1580 21023
rect 130 20907 1580 20937
rect 130 20821 1580 20851
rect 130 20735 1580 20765
rect 130 20649 1580 20679
rect 130 20563 1580 20593
rect 130 20477 1580 20507
rect 130 20391 1580 20421
rect 130 20305 1580 20335
rect 130 20219 1580 20249
rect 130 20133 1580 20163
rect 130 20047 1580 20077
rect 130 19961 1580 19991
rect 130 19875 1580 19905
rect 130 19789 1580 19819
rect 130 19703 1580 19733
rect 130 19617 1580 19647
rect 130 19531 1580 19561
rect 130 19445 1580 19475
rect 130 19359 1580 19389
rect 130 19273 1580 19303
rect 130 19187 1580 19217
rect 130 19101 1580 19131
rect 130 19015 1580 19045
rect 130 18929 1580 18959
rect 130 18843 1580 18873
rect 130 18757 1580 18787
rect 130 18671 1580 18701
rect 130 18585 1580 18615
rect 130 18499 1580 18529
rect 130 18413 1580 18443
rect 130 18327 1580 18357
rect 130 18241 1580 18271
rect 130 18155 1580 18185
rect 130 18069 1580 18099
rect 130 17983 1580 18013
rect 130 17897 1580 17927
rect 130 17811 1580 17841
rect 130 17725 1580 17755
rect 130 17639 1580 17669
rect 130 17553 1580 17583
rect 130 17467 1580 17497
rect 130 17381 1580 17411
rect 130 17295 1580 17325
rect 130 17209 1580 17239
rect 130 17123 1580 17153
rect 130 17037 1580 17067
rect 130 16951 1580 16981
rect 130 16865 1580 16895
rect 130 16779 1580 16809
rect 130 16693 1580 16723
rect 130 16607 1580 16637
rect 130 16521 1580 16551
rect 130 16435 1580 16465
rect 130 16349 1580 16379
rect 130 16263 1580 16293
rect 130 16177 1580 16207
rect 130 16091 1580 16121
rect 130 16005 1580 16035
rect 130 15919 1580 15949
rect 130 15833 1580 15863
rect 130 15747 1580 15777
rect 130 15661 1580 15691
rect 130 15575 1580 15605
rect 130 15489 1580 15519
rect 130 15403 1580 15433
rect 130 15317 1580 15347
rect 130 15231 1580 15261
rect 130 15145 1580 15175
rect 130 15059 1580 15089
rect 130 14973 1580 15003
rect 130 14887 1580 14917
rect 130 14801 1580 14831
rect 130 14715 1580 14745
rect 130 14629 1580 14659
rect 130 14543 1580 14573
rect 130 14457 1580 14487
rect 130 14371 1580 14401
rect 130 14285 1580 14315
rect 130 14199 1580 14229
rect 130 14113 1580 14143
rect 130 14027 1580 14057
rect 130 13941 1580 13971
rect 130 13855 1580 13885
rect 130 13769 1580 13799
rect 130 13683 1580 13713
rect 130 13597 1580 13627
rect 130 13511 1580 13541
rect 130 13425 1580 13455
rect 130 13339 1580 13369
rect 130 13253 1580 13283
rect 130 13167 1580 13197
rect 130 13081 1580 13111
rect 130 12995 1580 13025
rect 130 12909 1580 12939
rect 130 12823 1580 12853
rect 130 12737 1580 12767
rect 130 12651 1580 12681
rect 130 12565 1580 12595
rect 130 12479 1580 12509
rect 130 12393 1580 12423
rect 130 12307 1580 12337
rect 130 12221 1580 12251
rect 130 12135 1580 12165
rect 130 12049 1580 12079
rect 130 11963 1580 11993
rect 130 11877 1580 11907
rect 130 11791 1580 11821
rect 130 11705 1580 11735
rect 130 11619 1580 11649
rect 130 11533 1580 11563
rect 130 11447 1580 11477
rect 130 11361 1580 11391
rect 130 11275 1580 11305
rect 130 11189 1580 11219
rect 130 11103 1580 11133
rect 130 11017 1580 11047
rect 130 10931 1580 10961
rect 130 10845 1580 10875
rect 130 10759 1580 10789
rect 130 10673 1580 10703
rect 130 10587 1580 10617
rect 130 10501 1580 10531
rect 130 10415 1580 10445
rect 130 10329 1580 10359
rect 130 10243 1580 10273
rect 130 10157 1580 10187
rect 130 10071 1580 10101
rect 130 9985 1580 10015
rect 130 9899 1580 9929
rect 130 9813 1580 9843
rect 130 9727 1580 9757
rect 130 9641 1580 9671
rect 130 9555 1580 9585
rect 130 9469 1580 9499
rect 130 9383 1580 9413
rect 130 9297 1580 9327
rect 130 9211 1580 9241
rect 130 9125 1580 9155
rect 130 9039 1580 9069
rect 130 8953 1580 8983
rect 130 8867 1580 8897
rect 130 8781 1580 8811
rect 130 8695 1580 8725
rect 130 8609 1580 8639
rect 130 8523 1580 8553
rect 130 8437 1580 8467
rect 130 8351 1580 8381
rect 130 8265 1580 8295
rect 130 8179 1580 8209
rect 130 8093 1580 8123
rect 130 8007 1580 8037
rect 130 7921 1580 7951
rect 130 7835 1580 7865
rect 130 7749 1580 7779
rect 130 7663 1580 7693
rect 130 7577 1580 7607
rect 130 7491 1580 7521
rect 130 7405 1580 7435
rect 130 7319 1580 7349
rect 130 7233 1580 7263
rect 130 7147 1580 7177
rect 130 7061 1580 7091
rect 130 6975 1580 7005
rect 130 6889 1580 6919
rect 130 6803 1580 6833
rect 130 6717 1580 6747
rect 130 6631 1580 6661
rect 130 6545 1580 6575
rect 130 6459 1580 6489
rect 130 6373 1580 6403
rect 130 6287 1580 6317
rect 130 6201 1580 6231
rect 130 6115 1580 6145
rect 130 6029 1580 6059
rect 130 5943 1580 5973
rect 130 5857 1580 5887
rect 130 5771 1580 5801
rect 130 5685 1580 5715
rect 130 5599 1580 5629
rect 130 5513 1580 5543
rect 130 5427 1580 5457
rect 130 5341 1580 5371
rect 130 5255 1580 5285
rect 130 5169 1580 5199
rect 130 5083 1580 5113
rect 130 4997 1580 5027
rect 130 4911 1580 4941
rect 130 4825 1580 4855
rect 130 4739 1580 4769
rect 130 4653 1580 4683
rect 130 4567 1580 4597
rect 130 4481 1580 4511
rect 130 4395 1580 4425
rect 130 4309 1580 4339
rect 130 4223 1580 4253
rect 130 4137 1580 4167
rect 130 4051 1580 4081
rect 130 3965 1580 3995
rect 130 3879 1580 3909
rect 130 3793 1580 3823
rect 130 3707 1580 3737
rect 130 3621 1580 3651
rect 130 3535 1580 3565
rect 130 3449 1580 3479
rect 130 3363 1580 3393
rect 130 3277 1580 3307
rect 130 3191 1580 3221
rect 130 3105 1580 3135
rect 130 3019 1580 3049
rect 130 2933 1580 2963
rect 130 2847 1580 2877
rect 130 2761 1580 2791
rect 130 2675 1580 2705
rect 130 2589 1580 2619
rect 130 2503 1580 2533
rect 130 2417 1580 2447
rect 130 2331 1580 2361
rect 130 2245 1580 2275
rect 130 2159 1580 2189
rect 130 2073 1580 2103
rect 130 1987 1580 2017
rect 130 1901 1580 1931
rect 130 1815 1580 1845
rect 130 1729 1580 1759
rect 130 1643 1580 1673
rect 130 1557 1580 1587
rect 130 1471 1580 1501
rect 130 1385 1580 1415
rect 130 1299 1580 1329
rect 130 1213 1580 1243
rect 130 1127 1580 1157
rect 130 1041 1580 1071
rect 130 955 1580 985
rect 130 869 1580 899
rect 130 783 1580 813
rect 130 697 1580 727
rect 130 611 1580 641
rect 130 525 1580 555
rect 130 439 1580 469
rect 130 353 1580 383
rect 130 267 1580 297
rect 130 181 1580 211
<< pdiff >>
rect 130 43858 1580 43870
rect 130 43824 138 43858
rect 1572 43824 1580 43858
rect 130 43813 1580 43824
rect 130 43772 1580 43783
rect 130 43738 138 43772
rect 1572 43738 1580 43772
rect 130 43727 1580 43738
rect 130 43686 1580 43697
rect 130 43652 138 43686
rect 1572 43652 1580 43686
rect 130 43641 1580 43652
rect 130 43600 1580 43611
rect 130 43566 138 43600
rect 1572 43566 1580 43600
rect 130 43555 1580 43566
rect 130 43514 1580 43525
rect 130 43480 138 43514
rect 1572 43480 1580 43514
rect 130 43469 1580 43480
rect 130 43428 1580 43439
rect 130 43394 138 43428
rect 1572 43394 1580 43428
rect 130 43383 1580 43394
rect 130 43342 1580 43353
rect 130 43308 138 43342
rect 1572 43308 1580 43342
rect 130 43297 1580 43308
rect 130 43256 1580 43267
rect 130 43222 138 43256
rect 1572 43222 1580 43256
rect 130 43211 1580 43222
rect 130 43170 1580 43181
rect 130 43136 138 43170
rect 1572 43136 1580 43170
rect 130 43125 1580 43136
rect 130 43084 1580 43095
rect 130 43050 138 43084
rect 1572 43050 1580 43084
rect 130 43039 1580 43050
rect 130 42998 1580 43009
rect 130 42964 138 42998
rect 1572 42964 1580 42998
rect 130 42953 1580 42964
rect 130 42912 1580 42923
rect 130 42878 138 42912
rect 1572 42878 1580 42912
rect 130 42867 1580 42878
rect 130 42826 1580 42837
rect 130 42792 138 42826
rect 1572 42792 1580 42826
rect 130 42781 1580 42792
rect 130 42740 1580 42751
rect 130 42706 138 42740
rect 1572 42706 1580 42740
rect 130 42695 1580 42706
rect 130 42654 1580 42665
rect 130 42620 138 42654
rect 1572 42620 1580 42654
rect 130 42609 1580 42620
rect 130 42568 1580 42579
rect 130 42534 138 42568
rect 1572 42534 1580 42568
rect 130 42523 1580 42534
rect 130 42482 1580 42493
rect 130 42448 138 42482
rect 1572 42448 1580 42482
rect 130 42437 1580 42448
rect 130 42396 1580 42407
rect 130 42362 138 42396
rect 1572 42362 1580 42396
rect 130 42351 1580 42362
rect 130 42310 1580 42321
rect 130 42276 138 42310
rect 1572 42276 1580 42310
rect 130 42265 1580 42276
rect 130 42224 1580 42235
rect 130 42190 138 42224
rect 1572 42190 1580 42224
rect 130 42179 1580 42190
rect 130 42138 1580 42149
rect 130 42104 138 42138
rect 1572 42104 1580 42138
rect 130 42093 1580 42104
rect 130 42052 1580 42063
rect 130 42018 138 42052
rect 1572 42018 1580 42052
rect 130 42007 1580 42018
rect 130 41966 1580 41977
rect 130 41932 138 41966
rect 1572 41932 1580 41966
rect 130 41921 1580 41932
rect 130 41880 1580 41891
rect 130 41846 138 41880
rect 1572 41846 1580 41880
rect 130 41835 1580 41846
rect 130 41794 1580 41805
rect 130 41760 138 41794
rect 1572 41760 1580 41794
rect 130 41749 1580 41760
rect 130 41708 1580 41719
rect 130 41674 138 41708
rect 1572 41674 1580 41708
rect 130 41663 1580 41674
rect 130 41622 1580 41633
rect 130 41588 138 41622
rect 1572 41588 1580 41622
rect 130 41577 1580 41588
rect 130 41536 1580 41547
rect 130 41502 138 41536
rect 1572 41502 1580 41536
rect 130 41491 1580 41502
rect 130 41450 1580 41461
rect 130 41416 138 41450
rect 1572 41416 1580 41450
rect 130 41405 1580 41416
rect 130 41364 1580 41375
rect 130 41330 138 41364
rect 1572 41330 1580 41364
rect 130 41319 1580 41330
rect 130 41278 1580 41289
rect 130 41244 138 41278
rect 1572 41244 1580 41278
rect 130 41233 1580 41244
rect 130 41192 1580 41203
rect 130 41158 138 41192
rect 1572 41158 1580 41192
rect 130 41147 1580 41158
rect 130 41106 1580 41117
rect 130 41072 138 41106
rect 1572 41072 1580 41106
rect 130 41061 1580 41072
rect 130 41020 1580 41031
rect 130 40986 138 41020
rect 1572 40986 1580 41020
rect 130 40975 1580 40986
rect 130 40934 1580 40945
rect 130 40900 138 40934
rect 1572 40900 1580 40934
rect 130 40889 1580 40900
rect 130 40848 1580 40859
rect 130 40814 138 40848
rect 1572 40814 1580 40848
rect 130 40803 1580 40814
rect 130 40762 1580 40773
rect 130 40728 138 40762
rect 1572 40728 1580 40762
rect 130 40717 1580 40728
rect 130 40676 1580 40687
rect 130 40642 138 40676
rect 1572 40642 1580 40676
rect 130 40631 1580 40642
rect 130 40590 1580 40601
rect 130 40556 138 40590
rect 1572 40556 1580 40590
rect 130 40545 1580 40556
rect 130 40504 1580 40515
rect 130 40470 138 40504
rect 1572 40470 1580 40504
rect 130 40459 1580 40470
rect 130 40418 1580 40429
rect 130 40384 138 40418
rect 1572 40384 1580 40418
rect 130 40373 1580 40384
rect 130 40332 1580 40343
rect 130 40298 138 40332
rect 1572 40298 1580 40332
rect 130 40287 1580 40298
rect 130 40246 1580 40257
rect 130 40212 138 40246
rect 1572 40212 1580 40246
rect 130 40201 1580 40212
rect 130 40160 1580 40171
rect 130 40126 138 40160
rect 1572 40126 1580 40160
rect 130 40115 1580 40126
rect 130 40074 1580 40085
rect 130 40040 138 40074
rect 1572 40040 1580 40074
rect 130 40029 1580 40040
rect 130 39988 1580 39999
rect 130 39954 138 39988
rect 1572 39954 1580 39988
rect 130 39943 1580 39954
rect 130 39902 1580 39913
rect 130 39868 138 39902
rect 1572 39868 1580 39902
rect 130 39857 1580 39868
rect 130 39816 1580 39827
rect 130 39782 138 39816
rect 1572 39782 1580 39816
rect 130 39771 1580 39782
rect 130 39730 1580 39741
rect 130 39696 138 39730
rect 1572 39696 1580 39730
rect 130 39685 1580 39696
rect 130 39644 1580 39655
rect 130 39610 138 39644
rect 1572 39610 1580 39644
rect 130 39599 1580 39610
rect 130 39558 1580 39569
rect 130 39524 138 39558
rect 1572 39524 1580 39558
rect 130 39513 1580 39524
rect 130 39472 1580 39483
rect 130 39438 138 39472
rect 1572 39438 1580 39472
rect 130 39427 1580 39438
rect 130 39386 1580 39397
rect 130 39352 138 39386
rect 1572 39352 1580 39386
rect 130 39341 1580 39352
rect 130 39300 1580 39311
rect 130 39266 138 39300
rect 1572 39266 1580 39300
rect 130 39255 1580 39266
rect 130 39214 1580 39225
rect 130 39180 138 39214
rect 1572 39180 1580 39214
rect 130 39169 1580 39180
rect 130 39128 1580 39139
rect 130 39094 138 39128
rect 1572 39094 1580 39128
rect 130 39083 1580 39094
rect 130 39042 1580 39053
rect 130 39008 138 39042
rect 1572 39008 1580 39042
rect 130 38997 1580 39008
rect 130 38956 1580 38967
rect 130 38922 138 38956
rect 1572 38922 1580 38956
rect 130 38911 1580 38922
rect 130 38870 1580 38881
rect 130 38836 138 38870
rect 1572 38836 1580 38870
rect 130 38825 1580 38836
rect 130 38784 1580 38795
rect 130 38750 138 38784
rect 1572 38750 1580 38784
rect 130 38739 1580 38750
rect 130 38698 1580 38709
rect 130 38664 138 38698
rect 1572 38664 1580 38698
rect 130 38653 1580 38664
rect 130 38612 1580 38623
rect 130 38578 138 38612
rect 1572 38578 1580 38612
rect 130 38567 1580 38578
rect 130 38526 1580 38537
rect 130 38492 138 38526
rect 1572 38492 1580 38526
rect 130 38481 1580 38492
rect 130 38440 1580 38451
rect 130 38406 138 38440
rect 1572 38406 1580 38440
rect 130 38395 1580 38406
rect 130 38354 1580 38365
rect 130 38320 138 38354
rect 1572 38320 1580 38354
rect 130 38309 1580 38320
rect 130 38268 1580 38279
rect 130 38234 138 38268
rect 1572 38234 1580 38268
rect 130 38223 1580 38234
rect 130 38182 1580 38193
rect 130 38148 138 38182
rect 1572 38148 1580 38182
rect 130 38137 1580 38148
rect 130 38096 1580 38107
rect 130 38062 138 38096
rect 1572 38062 1580 38096
rect 130 38051 1580 38062
rect 130 38010 1580 38021
rect 130 37976 138 38010
rect 1572 37976 1580 38010
rect 130 37965 1580 37976
rect 130 37924 1580 37935
rect 130 37890 138 37924
rect 1572 37890 1580 37924
rect 130 37879 1580 37890
rect 130 37838 1580 37849
rect 130 37804 138 37838
rect 1572 37804 1580 37838
rect 130 37793 1580 37804
rect 130 37752 1580 37763
rect 130 37718 138 37752
rect 1572 37718 1580 37752
rect 130 37707 1580 37718
rect 130 37666 1580 37677
rect 130 37632 138 37666
rect 1572 37632 1580 37666
rect 130 37621 1580 37632
rect 130 37580 1580 37591
rect 130 37546 138 37580
rect 1572 37546 1580 37580
rect 130 37535 1580 37546
rect 130 37494 1580 37505
rect 130 37460 138 37494
rect 1572 37460 1580 37494
rect 130 37449 1580 37460
rect 130 37408 1580 37419
rect 130 37374 138 37408
rect 1572 37374 1580 37408
rect 130 37363 1580 37374
rect 130 37322 1580 37333
rect 130 37288 138 37322
rect 1572 37288 1580 37322
rect 130 37277 1580 37288
rect 130 37236 1580 37247
rect 130 37202 138 37236
rect 1572 37202 1580 37236
rect 130 37191 1580 37202
rect 130 37150 1580 37161
rect 130 37116 138 37150
rect 1572 37116 1580 37150
rect 130 37105 1580 37116
rect 130 37064 1580 37075
rect 130 37030 138 37064
rect 1572 37030 1580 37064
rect 130 37019 1580 37030
rect 130 36978 1580 36989
rect 130 36944 138 36978
rect 1572 36944 1580 36978
rect 130 36933 1580 36944
rect 130 36892 1580 36903
rect 130 36858 138 36892
rect 1572 36858 1580 36892
rect 130 36847 1580 36858
rect 130 36806 1580 36817
rect 130 36772 138 36806
rect 1572 36772 1580 36806
rect 130 36761 1580 36772
rect 130 36720 1580 36731
rect 130 36686 138 36720
rect 1572 36686 1580 36720
rect 130 36675 1580 36686
rect 130 36634 1580 36645
rect 130 36600 138 36634
rect 1572 36600 1580 36634
rect 130 36589 1580 36600
rect 130 36548 1580 36559
rect 130 36514 138 36548
rect 1572 36514 1580 36548
rect 130 36503 1580 36514
rect 130 36462 1580 36473
rect 130 36428 138 36462
rect 1572 36428 1580 36462
rect 130 36417 1580 36428
rect 130 36376 1580 36387
rect 130 36342 138 36376
rect 1572 36342 1580 36376
rect 130 36331 1580 36342
rect 130 36290 1580 36301
rect 130 36256 138 36290
rect 1572 36256 1580 36290
rect 130 36245 1580 36256
rect 130 36204 1580 36215
rect 130 36170 138 36204
rect 1572 36170 1580 36204
rect 130 36159 1580 36170
rect 130 36118 1580 36129
rect 130 36084 138 36118
rect 1572 36084 1580 36118
rect 130 36073 1580 36084
rect 130 36032 1580 36043
rect 130 35998 138 36032
rect 1572 35998 1580 36032
rect 130 35987 1580 35998
rect 130 35946 1580 35957
rect 130 35912 138 35946
rect 1572 35912 1580 35946
rect 130 35901 1580 35912
rect 130 35860 1580 35871
rect 130 35826 138 35860
rect 1572 35826 1580 35860
rect 130 35815 1580 35826
rect 130 35774 1580 35785
rect 130 35740 138 35774
rect 1572 35740 1580 35774
rect 130 35729 1580 35740
rect 130 35688 1580 35699
rect 130 35654 138 35688
rect 1572 35654 1580 35688
rect 130 35643 1580 35654
rect 130 35602 1580 35613
rect 130 35568 138 35602
rect 1572 35568 1580 35602
rect 130 35557 1580 35568
rect 130 35516 1580 35527
rect 130 35482 138 35516
rect 1572 35482 1580 35516
rect 130 35471 1580 35482
rect 130 35430 1580 35441
rect 130 35396 138 35430
rect 1572 35396 1580 35430
rect 130 35385 1580 35396
rect 130 35344 1580 35355
rect 130 35310 138 35344
rect 1572 35310 1580 35344
rect 130 35299 1580 35310
rect 130 35258 1580 35269
rect 130 35224 138 35258
rect 1572 35224 1580 35258
rect 130 35213 1580 35224
rect 130 35172 1580 35183
rect 130 35138 138 35172
rect 1572 35138 1580 35172
rect 130 35127 1580 35138
rect 130 35086 1580 35097
rect 130 35052 138 35086
rect 1572 35052 1580 35086
rect 130 35041 1580 35052
rect 130 35000 1580 35011
rect 130 34966 138 35000
rect 1572 34966 1580 35000
rect 130 34955 1580 34966
rect 130 34914 1580 34925
rect 130 34880 138 34914
rect 1572 34880 1580 34914
rect 130 34869 1580 34880
rect 130 34828 1580 34839
rect 130 34794 138 34828
rect 1572 34794 1580 34828
rect 130 34783 1580 34794
rect 130 34742 1580 34753
rect 130 34708 138 34742
rect 1572 34708 1580 34742
rect 130 34697 1580 34708
rect 130 34656 1580 34667
rect 130 34622 138 34656
rect 1572 34622 1580 34656
rect 130 34611 1580 34622
rect 130 34570 1580 34581
rect 130 34536 138 34570
rect 1572 34536 1580 34570
rect 130 34525 1580 34536
rect 130 34484 1580 34495
rect 130 34450 138 34484
rect 1572 34450 1580 34484
rect 130 34439 1580 34450
rect 130 34398 1580 34409
rect 130 34364 138 34398
rect 1572 34364 1580 34398
rect 130 34353 1580 34364
rect 130 34312 1580 34323
rect 130 34278 138 34312
rect 1572 34278 1580 34312
rect 130 34267 1580 34278
rect 130 34226 1580 34237
rect 130 34192 138 34226
rect 1572 34192 1580 34226
rect 130 34181 1580 34192
rect 130 34140 1580 34151
rect 130 34106 138 34140
rect 1572 34106 1580 34140
rect 130 34095 1580 34106
rect 130 34054 1580 34065
rect 130 34020 138 34054
rect 1572 34020 1580 34054
rect 130 34009 1580 34020
rect 130 33968 1580 33979
rect 130 33934 138 33968
rect 1572 33934 1580 33968
rect 130 33923 1580 33934
rect 130 33882 1580 33893
rect 130 33848 138 33882
rect 1572 33848 1580 33882
rect 130 33837 1580 33848
rect 130 33796 1580 33807
rect 130 33762 138 33796
rect 1572 33762 1580 33796
rect 130 33751 1580 33762
rect 130 33710 1580 33721
rect 130 33676 138 33710
rect 1572 33676 1580 33710
rect 130 33665 1580 33676
rect 130 33624 1580 33635
rect 130 33590 138 33624
rect 1572 33590 1580 33624
rect 130 33579 1580 33590
rect 130 33538 1580 33549
rect 130 33504 138 33538
rect 1572 33504 1580 33538
rect 130 33493 1580 33504
rect 130 33452 1580 33463
rect 130 33418 138 33452
rect 1572 33418 1580 33452
rect 130 33407 1580 33418
rect 130 33366 1580 33377
rect 130 33332 138 33366
rect 1572 33332 1580 33366
rect 130 33321 1580 33332
rect 130 33280 1580 33291
rect 130 33246 138 33280
rect 1572 33246 1580 33280
rect 130 33235 1580 33246
rect 130 33194 1580 33205
rect 130 33160 138 33194
rect 1572 33160 1580 33194
rect 130 33149 1580 33160
rect 130 33108 1580 33119
rect 130 33074 138 33108
rect 1572 33074 1580 33108
rect 130 33063 1580 33074
rect 130 33022 1580 33033
rect 130 32988 138 33022
rect 1572 32988 1580 33022
rect 130 32977 1580 32988
rect 130 32936 1580 32947
rect 130 32902 138 32936
rect 1572 32902 1580 32936
rect 130 32891 1580 32902
rect 130 32850 1580 32861
rect 130 32816 138 32850
rect 1572 32816 1580 32850
rect 130 32805 1580 32816
rect 130 32764 1580 32775
rect 130 32730 138 32764
rect 1572 32730 1580 32764
rect 130 32719 1580 32730
rect 130 32678 1580 32689
rect 130 32644 138 32678
rect 1572 32644 1580 32678
rect 130 32633 1580 32644
rect 130 32592 1580 32603
rect 130 32558 138 32592
rect 1572 32558 1580 32592
rect 130 32547 1580 32558
rect 130 32506 1580 32517
rect 130 32472 138 32506
rect 1572 32472 1580 32506
rect 130 32461 1580 32472
rect 130 32420 1580 32431
rect 130 32386 138 32420
rect 1572 32386 1580 32420
rect 130 32375 1580 32386
rect 130 32334 1580 32345
rect 130 32300 138 32334
rect 1572 32300 1580 32334
rect 130 32289 1580 32300
rect 130 32248 1580 32259
rect 130 32214 138 32248
rect 1572 32214 1580 32248
rect 130 32203 1580 32214
rect 130 32162 1580 32173
rect 130 32128 138 32162
rect 1572 32128 1580 32162
rect 130 32117 1580 32128
rect 130 32076 1580 32087
rect 130 32042 138 32076
rect 1572 32042 1580 32076
rect 130 32031 1580 32042
rect 130 31990 1580 32001
rect 130 31956 138 31990
rect 1572 31956 1580 31990
rect 130 31945 1580 31956
rect 130 31904 1580 31915
rect 130 31870 138 31904
rect 1572 31870 1580 31904
rect 130 31859 1580 31870
rect 130 31818 1580 31829
rect 130 31784 138 31818
rect 1572 31784 1580 31818
rect 130 31773 1580 31784
rect 130 31732 1580 31743
rect 130 31698 138 31732
rect 1572 31698 1580 31732
rect 130 31687 1580 31698
rect 130 31646 1580 31657
rect 130 31612 138 31646
rect 1572 31612 1580 31646
rect 130 31601 1580 31612
rect 130 31560 1580 31571
rect 130 31526 138 31560
rect 1572 31526 1580 31560
rect 130 31515 1580 31526
rect 130 31474 1580 31485
rect 130 31440 138 31474
rect 1572 31440 1580 31474
rect 130 31429 1580 31440
rect 130 31388 1580 31399
rect 130 31354 138 31388
rect 1572 31354 1580 31388
rect 130 31343 1580 31354
rect 130 31302 1580 31313
rect 130 31268 138 31302
rect 1572 31268 1580 31302
rect 130 31257 1580 31268
rect 130 31216 1580 31227
rect 130 31182 138 31216
rect 1572 31182 1580 31216
rect 130 31171 1580 31182
rect 130 31130 1580 31141
rect 130 31096 138 31130
rect 1572 31096 1580 31130
rect 130 31085 1580 31096
rect 130 31044 1580 31055
rect 130 31010 138 31044
rect 1572 31010 1580 31044
rect 130 30999 1580 31010
rect 130 30958 1580 30969
rect 130 30924 138 30958
rect 1572 30924 1580 30958
rect 130 30913 1580 30924
rect 130 30872 1580 30883
rect 130 30838 138 30872
rect 1572 30838 1580 30872
rect 130 30827 1580 30838
rect 130 30786 1580 30797
rect 130 30752 138 30786
rect 1572 30752 1580 30786
rect 130 30741 1580 30752
rect 130 30700 1580 30711
rect 130 30666 138 30700
rect 1572 30666 1580 30700
rect 130 30655 1580 30666
rect 130 30614 1580 30625
rect 130 30580 138 30614
rect 1572 30580 1580 30614
rect 130 30569 1580 30580
rect 130 30528 1580 30539
rect 130 30494 138 30528
rect 1572 30494 1580 30528
rect 130 30483 1580 30494
rect 130 30442 1580 30453
rect 130 30408 138 30442
rect 1572 30408 1580 30442
rect 130 30397 1580 30408
rect 130 30356 1580 30367
rect 130 30322 138 30356
rect 1572 30322 1580 30356
rect 130 30311 1580 30322
rect 130 30270 1580 30281
rect 130 30236 138 30270
rect 1572 30236 1580 30270
rect 130 30225 1580 30236
rect 130 30184 1580 30195
rect 130 30150 138 30184
rect 1572 30150 1580 30184
rect 130 30139 1580 30150
rect 130 30098 1580 30109
rect 130 30064 138 30098
rect 1572 30064 1580 30098
rect 130 30053 1580 30064
rect 130 30012 1580 30023
rect 130 29978 138 30012
rect 1572 29978 1580 30012
rect 130 29967 1580 29978
rect 130 29926 1580 29937
rect 130 29892 138 29926
rect 1572 29892 1580 29926
rect 130 29881 1580 29892
rect 130 29840 1580 29851
rect 130 29806 138 29840
rect 1572 29806 1580 29840
rect 130 29795 1580 29806
rect 130 29754 1580 29765
rect 130 29720 138 29754
rect 1572 29720 1580 29754
rect 130 29709 1580 29720
rect 130 29668 1580 29679
rect 130 29634 138 29668
rect 1572 29634 1580 29668
rect 130 29623 1580 29634
rect 130 29582 1580 29593
rect 130 29548 138 29582
rect 1572 29548 1580 29582
rect 130 29537 1580 29548
rect 130 29496 1580 29507
rect 130 29462 138 29496
rect 1572 29462 1580 29496
rect 130 29451 1580 29462
rect 130 29410 1580 29421
rect 130 29376 138 29410
rect 1572 29376 1580 29410
rect 130 29365 1580 29376
rect 130 29324 1580 29335
rect 130 29290 138 29324
rect 1572 29290 1580 29324
rect 130 29279 1580 29290
rect 130 29238 1580 29249
rect 130 29204 138 29238
rect 1572 29204 1580 29238
rect 130 29193 1580 29204
rect 130 29152 1580 29163
rect 130 29118 138 29152
rect 1572 29118 1580 29152
rect 130 29107 1580 29118
rect 130 29066 1580 29077
rect 130 29032 138 29066
rect 1572 29032 1580 29066
rect 130 29021 1580 29032
rect 130 28980 1580 28991
rect 130 28946 138 28980
rect 1572 28946 1580 28980
rect 130 28935 1580 28946
rect 130 28894 1580 28905
rect 130 28860 138 28894
rect 1572 28860 1580 28894
rect 130 28849 1580 28860
rect 130 28808 1580 28819
rect 130 28774 138 28808
rect 1572 28774 1580 28808
rect 130 28763 1580 28774
rect 130 28722 1580 28733
rect 130 28688 138 28722
rect 1572 28688 1580 28722
rect 130 28677 1580 28688
rect 130 28636 1580 28647
rect 130 28602 138 28636
rect 1572 28602 1580 28636
rect 130 28591 1580 28602
rect 130 28550 1580 28561
rect 130 28516 138 28550
rect 1572 28516 1580 28550
rect 130 28505 1580 28516
rect 130 28464 1580 28475
rect 130 28430 138 28464
rect 1572 28430 1580 28464
rect 130 28419 1580 28430
rect 130 28378 1580 28389
rect 130 28344 138 28378
rect 1572 28344 1580 28378
rect 130 28333 1580 28344
rect 130 28292 1580 28303
rect 130 28258 138 28292
rect 1572 28258 1580 28292
rect 130 28247 1580 28258
rect 130 28206 1580 28217
rect 130 28172 138 28206
rect 1572 28172 1580 28206
rect 130 28161 1580 28172
rect 130 28120 1580 28131
rect 130 28086 138 28120
rect 1572 28086 1580 28120
rect 130 28075 1580 28086
rect 130 28034 1580 28045
rect 130 28000 138 28034
rect 1572 28000 1580 28034
rect 130 27989 1580 28000
rect 130 27948 1580 27959
rect 130 27914 138 27948
rect 1572 27914 1580 27948
rect 130 27903 1580 27914
rect 130 27862 1580 27873
rect 130 27828 138 27862
rect 1572 27828 1580 27862
rect 130 27817 1580 27828
rect 130 27776 1580 27787
rect 130 27742 138 27776
rect 1572 27742 1580 27776
rect 130 27731 1580 27742
rect 130 27690 1580 27701
rect 130 27656 138 27690
rect 1572 27656 1580 27690
rect 130 27645 1580 27656
rect 130 27604 1580 27615
rect 130 27570 138 27604
rect 1572 27570 1580 27604
rect 130 27559 1580 27570
rect 130 27518 1580 27529
rect 130 27484 138 27518
rect 1572 27484 1580 27518
rect 130 27473 1580 27484
rect 130 27432 1580 27443
rect 130 27398 138 27432
rect 1572 27398 1580 27432
rect 130 27387 1580 27398
rect 130 27346 1580 27357
rect 130 27312 138 27346
rect 1572 27312 1580 27346
rect 130 27301 1580 27312
rect 130 27260 1580 27271
rect 130 27226 138 27260
rect 1572 27226 1580 27260
rect 130 27215 1580 27226
rect 130 27174 1580 27185
rect 130 27140 138 27174
rect 1572 27140 1580 27174
rect 130 27129 1580 27140
rect 130 27088 1580 27099
rect 130 27054 138 27088
rect 1572 27054 1580 27088
rect 130 27043 1580 27054
rect 130 27002 1580 27013
rect 130 26968 138 27002
rect 1572 26968 1580 27002
rect 130 26957 1580 26968
rect 130 26916 1580 26927
rect 130 26882 138 26916
rect 1572 26882 1580 26916
rect 130 26871 1580 26882
rect 130 26830 1580 26841
rect 130 26796 138 26830
rect 1572 26796 1580 26830
rect 130 26785 1580 26796
rect 130 26744 1580 26755
rect 130 26710 138 26744
rect 1572 26710 1580 26744
rect 130 26699 1580 26710
rect 130 26658 1580 26669
rect 130 26624 138 26658
rect 1572 26624 1580 26658
rect 130 26613 1580 26624
rect 130 26572 1580 26583
rect 130 26538 138 26572
rect 1572 26538 1580 26572
rect 130 26527 1580 26538
rect 130 26486 1580 26497
rect 130 26452 138 26486
rect 1572 26452 1580 26486
rect 130 26441 1580 26452
rect 130 26400 1580 26411
rect 130 26366 138 26400
rect 1572 26366 1580 26400
rect 130 26355 1580 26366
rect 130 26314 1580 26325
rect 130 26280 138 26314
rect 1572 26280 1580 26314
rect 130 26269 1580 26280
rect 130 26228 1580 26239
rect 130 26194 138 26228
rect 1572 26194 1580 26228
rect 130 26183 1580 26194
rect 130 26142 1580 26153
rect 130 26108 138 26142
rect 1572 26108 1580 26142
rect 130 26097 1580 26108
rect 130 26056 1580 26067
rect 130 26022 138 26056
rect 1572 26022 1580 26056
rect 130 26011 1580 26022
rect 130 25970 1580 25981
rect 130 25936 138 25970
rect 1572 25936 1580 25970
rect 130 25925 1580 25936
rect 130 25884 1580 25895
rect 130 25850 138 25884
rect 1572 25850 1580 25884
rect 130 25839 1580 25850
rect 130 25798 1580 25809
rect 130 25764 138 25798
rect 1572 25764 1580 25798
rect 130 25753 1580 25764
rect 130 25712 1580 25723
rect 130 25678 138 25712
rect 1572 25678 1580 25712
rect 130 25667 1580 25678
rect 130 25626 1580 25637
rect 130 25592 138 25626
rect 1572 25592 1580 25626
rect 130 25581 1580 25592
rect 130 25540 1580 25551
rect 130 25506 138 25540
rect 1572 25506 1580 25540
rect 130 25495 1580 25506
rect 130 25454 1580 25465
rect 130 25420 138 25454
rect 1572 25420 1580 25454
rect 130 25409 1580 25420
rect 130 25368 1580 25379
rect 130 25334 138 25368
rect 1572 25334 1580 25368
rect 130 25323 1580 25334
rect 130 25282 1580 25293
rect 130 25248 138 25282
rect 1572 25248 1580 25282
rect 130 25237 1580 25248
rect 130 25196 1580 25207
rect 130 25162 138 25196
rect 1572 25162 1580 25196
rect 130 25151 1580 25162
rect 130 25110 1580 25121
rect 130 25076 138 25110
rect 1572 25076 1580 25110
rect 130 25065 1580 25076
rect 130 25024 1580 25035
rect 130 24990 138 25024
rect 1572 24990 1580 25024
rect 130 24979 1580 24990
rect 130 24938 1580 24949
rect 130 24904 138 24938
rect 1572 24904 1580 24938
rect 130 24893 1580 24904
rect 130 24852 1580 24863
rect 130 24818 138 24852
rect 1572 24818 1580 24852
rect 130 24807 1580 24818
rect 130 24766 1580 24777
rect 130 24732 138 24766
rect 1572 24732 1580 24766
rect 130 24721 1580 24732
rect 130 24680 1580 24691
rect 130 24646 138 24680
rect 1572 24646 1580 24680
rect 130 24635 1580 24646
rect 130 24594 1580 24605
rect 130 24560 138 24594
rect 1572 24560 1580 24594
rect 130 24549 1580 24560
rect 130 24508 1580 24519
rect 130 24474 138 24508
rect 1572 24474 1580 24508
rect 130 24463 1580 24474
rect 130 24422 1580 24433
rect 130 24388 138 24422
rect 1572 24388 1580 24422
rect 130 24377 1580 24388
rect 130 24336 1580 24347
rect 130 24302 138 24336
rect 1572 24302 1580 24336
rect 130 24291 1580 24302
rect 130 24250 1580 24261
rect 130 24216 138 24250
rect 1572 24216 1580 24250
rect 130 24205 1580 24216
rect 130 24164 1580 24175
rect 130 24130 138 24164
rect 1572 24130 1580 24164
rect 130 24119 1580 24130
rect 130 24078 1580 24089
rect 130 24044 138 24078
rect 1572 24044 1580 24078
rect 130 24033 1580 24044
rect 130 23992 1580 24003
rect 130 23958 138 23992
rect 1572 23958 1580 23992
rect 130 23947 1580 23958
rect 130 23906 1580 23917
rect 130 23872 138 23906
rect 1572 23872 1580 23906
rect 130 23861 1580 23872
rect 130 23820 1580 23831
rect 130 23786 138 23820
rect 1572 23786 1580 23820
rect 130 23775 1580 23786
rect 130 23734 1580 23745
rect 130 23700 138 23734
rect 1572 23700 1580 23734
rect 130 23689 1580 23700
rect 130 23648 1580 23659
rect 130 23614 138 23648
rect 1572 23614 1580 23648
rect 130 23603 1580 23614
rect 130 23562 1580 23573
rect 130 23528 138 23562
rect 1572 23528 1580 23562
rect 130 23517 1580 23528
rect 130 23476 1580 23487
rect 130 23442 138 23476
rect 1572 23442 1580 23476
rect 130 23431 1580 23442
rect 130 23390 1580 23401
rect 130 23356 138 23390
rect 1572 23356 1580 23390
rect 130 23345 1580 23356
rect 130 23304 1580 23315
rect 130 23270 138 23304
rect 1572 23270 1580 23304
rect 130 23259 1580 23270
rect 130 23218 1580 23229
rect 130 23184 138 23218
rect 1572 23184 1580 23218
rect 130 23173 1580 23184
rect 130 23132 1580 23143
rect 130 23098 138 23132
rect 1572 23098 1580 23132
rect 130 23087 1580 23098
rect 130 23046 1580 23057
rect 130 23012 138 23046
rect 1572 23012 1580 23046
rect 130 23001 1580 23012
rect 130 22960 1580 22971
rect 130 22926 138 22960
rect 1572 22926 1580 22960
rect 130 22915 1580 22926
rect 130 22874 1580 22885
rect 130 22840 138 22874
rect 1572 22840 1580 22874
rect 130 22829 1580 22840
rect 130 22788 1580 22799
rect 130 22754 138 22788
rect 1572 22754 1580 22788
rect 130 22743 1580 22754
rect 130 22702 1580 22713
rect 130 22668 138 22702
rect 1572 22668 1580 22702
rect 130 22657 1580 22668
rect 130 22616 1580 22627
rect 130 22582 138 22616
rect 1572 22582 1580 22616
rect 130 22571 1580 22582
rect 130 22530 1580 22541
rect 130 22496 138 22530
rect 1572 22496 1580 22530
rect 130 22485 1580 22496
rect 130 22444 1580 22455
rect 130 22410 138 22444
rect 1572 22410 1580 22444
rect 130 22399 1580 22410
rect 130 22358 1580 22369
rect 130 22324 138 22358
rect 1572 22324 1580 22358
rect 130 22313 1580 22324
rect 130 22272 1580 22283
rect 130 22238 138 22272
rect 1572 22238 1580 22272
rect 130 22227 1580 22238
rect 130 22186 1580 22197
rect 130 22152 138 22186
rect 1572 22152 1580 22186
rect 130 22141 1580 22152
rect 130 22100 1580 22111
rect 130 22066 138 22100
rect 1572 22066 1580 22100
rect 130 22055 1580 22066
rect 130 22014 1580 22025
rect 130 21980 138 22014
rect 1572 21980 1580 22014
rect 130 21969 1580 21980
rect 130 21928 1580 21939
rect 130 21894 138 21928
rect 1572 21894 1580 21928
rect 130 21883 1580 21894
rect 130 21842 1580 21853
rect 130 21808 138 21842
rect 1572 21808 1580 21842
rect 130 21797 1580 21808
rect 130 21756 1580 21767
rect 130 21722 138 21756
rect 1572 21722 1580 21756
rect 130 21711 1580 21722
rect 130 21670 1580 21681
rect 130 21636 138 21670
rect 1572 21636 1580 21670
rect 130 21625 1580 21636
rect 130 21584 1580 21595
rect 130 21550 138 21584
rect 1572 21550 1580 21584
rect 130 21539 1580 21550
rect 130 21498 1580 21509
rect 130 21464 138 21498
rect 1572 21464 1580 21498
rect 130 21453 1580 21464
rect 130 21412 1580 21423
rect 130 21378 138 21412
rect 1572 21378 1580 21412
rect 130 21367 1580 21378
rect 130 21326 1580 21337
rect 130 21292 138 21326
rect 1572 21292 1580 21326
rect 130 21281 1580 21292
rect 130 21240 1580 21251
rect 130 21206 138 21240
rect 1572 21206 1580 21240
rect 130 21195 1580 21206
rect 130 21154 1580 21165
rect 130 21120 138 21154
rect 1572 21120 1580 21154
rect 130 21109 1580 21120
rect 130 21068 1580 21079
rect 130 21034 138 21068
rect 1572 21034 1580 21068
rect 130 21023 1580 21034
rect 130 20982 1580 20993
rect 130 20948 138 20982
rect 1572 20948 1580 20982
rect 130 20937 1580 20948
rect 130 20896 1580 20907
rect 130 20862 138 20896
rect 1572 20862 1580 20896
rect 130 20851 1580 20862
rect 130 20810 1580 20821
rect 130 20776 138 20810
rect 1572 20776 1580 20810
rect 130 20765 1580 20776
rect 130 20724 1580 20735
rect 130 20690 138 20724
rect 1572 20690 1580 20724
rect 130 20679 1580 20690
rect 130 20638 1580 20649
rect 130 20604 138 20638
rect 1572 20604 1580 20638
rect 130 20593 1580 20604
rect 130 20552 1580 20563
rect 130 20518 138 20552
rect 1572 20518 1580 20552
rect 130 20507 1580 20518
rect 130 20466 1580 20477
rect 130 20432 138 20466
rect 1572 20432 1580 20466
rect 130 20421 1580 20432
rect 130 20380 1580 20391
rect 130 20346 138 20380
rect 1572 20346 1580 20380
rect 130 20335 1580 20346
rect 130 20294 1580 20305
rect 130 20260 138 20294
rect 1572 20260 1580 20294
rect 130 20249 1580 20260
rect 130 20208 1580 20219
rect 130 20174 138 20208
rect 1572 20174 1580 20208
rect 130 20163 1580 20174
rect 130 20122 1580 20133
rect 130 20088 138 20122
rect 1572 20088 1580 20122
rect 130 20077 1580 20088
rect 130 20036 1580 20047
rect 130 20002 138 20036
rect 1572 20002 1580 20036
rect 130 19991 1580 20002
rect 130 19950 1580 19961
rect 130 19916 138 19950
rect 1572 19916 1580 19950
rect 130 19905 1580 19916
rect 130 19864 1580 19875
rect 130 19830 138 19864
rect 1572 19830 1580 19864
rect 130 19819 1580 19830
rect 130 19778 1580 19789
rect 130 19744 138 19778
rect 1572 19744 1580 19778
rect 130 19733 1580 19744
rect 130 19692 1580 19703
rect 130 19658 138 19692
rect 1572 19658 1580 19692
rect 130 19647 1580 19658
rect 130 19606 1580 19617
rect 130 19572 138 19606
rect 1572 19572 1580 19606
rect 130 19561 1580 19572
rect 130 19520 1580 19531
rect 130 19486 138 19520
rect 1572 19486 1580 19520
rect 130 19475 1580 19486
rect 130 19434 1580 19445
rect 130 19400 138 19434
rect 1572 19400 1580 19434
rect 130 19389 1580 19400
rect 130 19348 1580 19359
rect 130 19314 138 19348
rect 1572 19314 1580 19348
rect 130 19303 1580 19314
rect 130 19262 1580 19273
rect 130 19228 138 19262
rect 1572 19228 1580 19262
rect 130 19217 1580 19228
rect 130 19176 1580 19187
rect 130 19142 138 19176
rect 1572 19142 1580 19176
rect 130 19131 1580 19142
rect 130 19090 1580 19101
rect 130 19056 138 19090
rect 1572 19056 1580 19090
rect 130 19045 1580 19056
rect 130 19004 1580 19015
rect 130 18970 138 19004
rect 1572 18970 1580 19004
rect 130 18959 1580 18970
rect 130 18918 1580 18929
rect 130 18884 138 18918
rect 1572 18884 1580 18918
rect 130 18873 1580 18884
rect 130 18832 1580 18843
rect 130 18798 138 18832
rect 1572 18798 1580 18832
rect 130 18787 1580 18798
rect 130 18746 1580 18757
rect 130 18712 138 18746
rect 1572 18712 1580 18746
rect 130 18701 1580 18712
rect 130 18660 1580 18671
rect 130 18626 138 18660
rect 1572 18626 1580 18660
rect 130 18615 1580 18626
rect 130 18574 1580 18585
rect 130 18540 138 18574
rect 1572 18540 1580 18574
rect 130 18529 1580 18540
rect 130 18488 1580 18499
rect 130 18454 138 18488
rect 1572 18454 1580 18488
rect 130 18443 1580 18454
rect 130 18402 1580 18413
rect 130 18368 138 18402
rect 1572 18368 1580 18402
rect 130 18357 1580 18368
rect 130 18316 1580 18327
rect 130 18282 138 18316
rect 1572 18282 1580 18316
rect 130 18271 1580 18282
rect 130 18230 1580 18241
rect 130 18196 138 18230
rect 1572 18196 1580 18230
rect 130 18185 1580 18196
rect 130 18144 1580 18155
rect 130 18110 138 18144
rect 1572 18110 1580 18144
rect 130 18099 1580 18110
rect 130 18058 1580 18069
rect 130 18024 138 18058
rect 1572 18024 1580 18058
rect 130 18013 1580 18024
rect 130 17972 1580 17983
rect 130 17938 138 17972
rect 1572 17938 1580 17972
rect 130 17927 1580 17938
rect 130 17886 1580 17897
rect 130 17852 138 17886
rect 1572 17852 1580 17886
rect 130 17841 1580 17852
rect 130 17800 1580 17811
rect 130 17766 138 17800
rect 1572 17766 1580 17800
rect 130 17755 1580 17766
rect 130 17714 1580 17725
rect 130 17680 138 17714
rect 1572 17680 1580 17714
rect 130 17669 1580 17680
rect 130 17628 1580 17639
rect 130 17594 138 17628
rect 1572 17594 1580 17628
rect 130 17583 1580 17594
rect 130 17542 1580 17553
rect 130 17508 138 17542
rect 1572 17508 1580 17542
rect 130 17497 1580 17508
rect 130 17456 1580 17467
rect 130 17422 138 17456
rect 1572 17422 1580 17456
rect 130 17411 1580 17422
rect 130 17370 1580 17381
rect 130 17336 138 17370
rect 1572 17336 1580 17370
rect 130 17325 1580 17336
rect 130 17284 1580 17295
rect 130 17250 138 17284
rect 1572 17250 1580 17284
rect 130 17239 1580 17250
rect 130 17198 1580 17209
rect 130 17164 138 17198
rect 1572 17164 1580 17198
rect 130 17153 1580 17164
rect 130 17112 1580 17123
rect 130 17078 138 17112
rect 1572 17078 1580 17112
rect 130 17067 1580 17078
rect 130 17026 1580 17037
rect 130 16992 138 17026
rect 1572 16992 1580 17026
rect 130 16981 1580 16992
rect 130 16940 1580 16951
rect 130 16906 138 16940
rect 1572 16906 1580 16940
rect 130 16895 1580 16906
rect 130 16854 1580 16865
rect 130 16820 138 16854
rect 1572 16820 1580 16854
rect 130 16809 1580 16820
rect 130 16768 1580 16779
rect 130 16734 138 16768
rect 1572 16734 1580 16768
rect 130 16723 1580 16734
rect 130 16682 1580 16693
rect 130 16648 138 16682
rect 1572 16648 1580 16682
rect 130 16637 1580 16648
rect 130 16596 1580 16607
rect 130 16562 138 16596
rect 1572 16562 1580 16596
rect 130 16551 1580 16562
rect 130 16510 1580 16521
rect 130 16476 138 16510
rect 1572 16476 1580 16510
rect 130 16465 1580 16476
rect 130 16424 1580 16435
rect 130 16390 138 16424
rect 1572 16390 1580 16424
rect 130 16379 1580 16390
rect 130 16338 1580 16349
rect 130 16304 138 16338
rect 1572 16304 1580 16338
rect 130 16293 1580 16304
rect 130 16252 1580 16263
rect 130 16218 138 16252
rect 1572 16218 1580 16252
rect 130 16207 1580 16218
rect 130 16166 1580 16177
rect 130 16132 138 16166
rect 1572 16132 1580 16166
rect 130 16121 1580 16132
rect 130 16080 1580 16091
rect 130 16046 138 16080
rect 1572 16046 1580 16080
rect 130 16035 1580 16046
rect 130 15994 1580 16005
rect 130 15960 138 15994
rect 1572 15960 1580 15994
rect 130 15949 1580 15960
rect 130 15908 1580 15919
rect 130 15874 138 15908
rect 1572 15874 1580 15908
rect 130 15863 1580 15874
rect 130 15822 1580 15833
rect 130 15788 138 15822
rect 1572 15788 1580 15822
rect 130 15777 1580 15788
rect 130 15736 1580 15747
rect 130 15702 138 15736
rect 1572 15702 1580 15736
rect 130 15691 1580 15702
rect 130 15650 1580 15661
rect 130 15616 138 15650
rect 1572 15616 1580 15650
rect 130 15605 1580 15616
rect 130 15564 1580 15575
rect 130 15530 138 15564
rect 1572 15530 1580 15564
rect 130 15519 1580 15530
rect 130 15478 1580 15489
rect 130 15444 138 15478
rect 1572 15444 1580 15478
rect 130 15433 1580 15444
rect 130 15392 1580 15403
rect 130 15358 138 15392
rect 1572 15358 1580 15392
rect 130 15347 1580 15358
rect 130 15306 1580 15317
rect 130 15272 138 15306
rect 1572 15272 1580 15306
rect 130 15261 1580 15272
rect 130 15220 1580 15231
rect 130 15186 138 15220
rect 1572 15186 1580 15220
rect 130 15175 1580 15186
rect 130 15134 1580 15145
rect 130 15100 138 15134
rect 1572 15100 1580 15134
rect 130 15089 1580 15100
rect 130 15048 1580 15059
rect 130 15014 138 15048
rect 1572 15014 1580 15048
rect 130 15003 1580 15014
rect 130 14962 1580 14973
rect 130 14928 138 14962
rect 1572 14928 1580 14962
rect 130 14917 1580 14928
rect 130 14876 1580 14887
rect 130 14842 138 14876
rect 1572 14842 1580 14876
rect 130 14831 1580 14842
rect 130 14790 1580 14801
rect 130 14756 138 14790
rect 1572 14756 1580 14790
rect 130 14745 1580 14756
rect 130 14704 1580 14715
rect 130 14670 138 14704
rect 1572 14670 1580 14704
rect 130 14659 1580 14670
rect 130 14618 1580 14629
rect 130 14584 138 14618
rect 1572 14584 1580 14618
rect 130 14573 1580 14584
rect 130 14532 1580 14543
rect 130 14498 138 14532
rect 1572 14498 1580 14532
rect 130 14487 1580 14498
rect 130 14446 1580 14457
rect 130 14412 138 14446
rect 1572 14412 1580 14446
rect 130 14401 1580 14412
rect 130 14360 1580 14371
rect 130 14326 138 14360
rect 1572 14326 1580 14360
rect 130 14315 1580 14326
rect 130 14274 1580 14285
rect 130 14240 138 14274
rect 1572 14240 1580 14274
rect 130 14229 1580 14240
rect 130 14188 1580 14199
rect 130 14154 138 14188
rect 1572 14154 1580 14188
rect 130 14143 1580 14154
rect 130 14102 1580 14113
rect 130 14068 138 14102
rect 1572 14068 1580 14102
rect 130 14057 1580 14068
rect 130 14016 1580 14027
rect 130 13982 138 14016
rect 1572 13982 1580 14016
rect 130 13971 1580 13982
rect 130 13930 1580 13941
rect 130 13896 138 13930
rect 1572 13896 1580 13930
rect 130 13885 1580 13896
rect 130 13844 1580 13855
rect 130 13810 138 13844
rect 1572 13810 1580 13844
rect 130 13799 1580 13810
rect 130 13758 1580 13769
rect 130 13724 138 13758
rect 1572 13724 1580 13758
rect 130 13713 1580 13724
rect 130 13672 1580 13683
rect 130 13638 138 13672
rect 1572 13638 1580 13672
rect 130 13627 1580 13638
rect 130 13586 1580 13597
rect 130 13552 138 13586
rect 1572 13552 1580 13586
rect 130 13541 1580 13552
rect 130 13500 1580 13511
rect 130 13466 138 13500
rect 1572 13466 1580 13500
rect 130 13455 1580 13466
rect 130 13414 1580 13425
rect 130 13380 138 13414
rect 1572 13380 1580 13414
rect 130 13369 1580 13380
rect 130 13328 1580 13339
rect 130 13294 138 13328
rect 1572 13294 1580 13328
rect 130 13283 1580 13294
rect 130 13242 1580 13253
rect 130 13208 138 13242
rect 1572 13208 1580 13242
rect 130 13197 1580 13208
rect 130 13156 1580 13167
rect 130 13122 138 13156
rect 1572 13122 1580 13156
rect 130 13111 1580 13122
rect 130 13070 1580 13081
rect 130 13036 138 13070
rect 1572 13036 1580 13070
rect 130 13025 1580 13036
rect 130 12984 1580 12995
rect 130 12950 138 12984
rect 1572 12950 1580 12984
rect 130 12939 1580 12950
rect 130 12898 1580 12909
rect 130 12864 138 12898
rect 1572 12864 1580 12898
rect 130 12853 1580 12864
rect 130 12812 1580 12823
rect 130 12778 138 12812
rect 1572 12778 1580 12812
rect 130 12767 1580 12778
rect 130 12726 1580 12737
rect 130 12692 138 12726
rect 1572 12692 1580 12726
rect 130 12681 1580 12692
rect 130 12640 1580 12651
rect 130 12606 138 12640
rect 1572 12606 1580 12640
rect 130 12595 1580 12606
rect 130 12554 1580 12565
rect 130 12520 138 12554
rect 1572 12520 1580 12554
rect 130 12509 1580 12520
rect 130 12468 1580 12479
rect 130 12434 138 12468
rect 1572 12434 1580 12468
rect 130 12423 1580 12434
rect 130 12382 1580 12393
rect 130 12348 138 12382
rect 1572 12348 1580 12382
rect 130 12337 1580 12348
rect 130 12296 1580 12307
rect 130 12262 138 12296
rect 1572 12262 1580 12296
rect 130 12251 1580 12262
rect 130 12210 1580 12221
rect 130 12176 138 12210
rect 1572 12176 1580 12210
rect 130 12165 1580 12176
rect 130 12124 1580 12135
rect 130 12090 138 12124
rect 1572 12090 1580 12124
rect 130 12079 1580 12090
rect 130 12038 1580 12049
rect 130 12004 138 12038
rect 1572 12004 1580 12038
rect 130 11993 1580 12004
rect 130 11952 1580 11963
rect 130 11918 138 11952
rect 1572 11918 1580 11952
rect 130 11907 1580 11918
rect 130 11866 1580 11877
rect 130 11832 138 11866
rect 1572 11832 1580 11866
rect 130 11821 1580 11832
rect 130 11780 1580 11791
rect 130 11746 138 11780
rect 1572 11746 1580 11780
rect 130 11735 1580 11746
rect 130 11694 1580 11705
rect 130 11660 138 11694
rect 1572 11660 1580 11694
rect 130 11649 1580 11660
rect 130 11608 1580 11619
rect 130 11574 138 11608
rect 1572 11574 1580 11608
rect 130 11563 1580 11574
rect 130 11522 1580 11533
rect 130 11488 138 11522
rect 1572 11488 1580 11522
rect 130 11477 1580 11488
rect 130 11436 1580 11447
rect 130 11402 138 11436
rect 1572 11402 1580 11436
rect 130 11391 1580 11402
rect 130 11350 1580 11361
rect 130 11316 138 11350
rect 1572 11316 1580 11350
rect 130 11305 1580 11316
rect 130 11264 1580 11275
rect 130 11230 138 11264
rect 1572 11230 1580 11264
rect 130 11219 1580 11230
rect 130 11178 1580 11189
rect 130 11144 138 11178
rect 1572 11144 1580 11178
rect 130 11133 1580 11144
rect 130 11092 1580 11103
rect 130 11058 138 11092
rect 1572 11058 1580 11092
rect 130 11047 1580 11058
rect 130 11006 1580 11017
rect 130 10972 138 11006
rect 1572 10972 1580 11006
rect 130 10961 1580 10972
rect 130 10920 1580 10931
rect 130 10886 138 10920
rect 1572 10886 1580 10920
rect 130 10875 1580 10886
rect 130 10834 1580 10845
rect 130 10800 138 10834
rect 1572 10800 1580 10834
rect 130 10789 1580 10800
rect 130 10748 1580 10759
rect 130 10714 138 10748
rect 1572 10714 1580 10748
rect 130 10703 1580 10714
rect 130 10662 1580 10673
rect 130 10628 138 10662
rect 1572 10628 1580 10662
rect 130 10617 1580 10628
rect 130 10576 1580 10587
rect 130 10542 138 10576
rect 1572 10542 1580 10576
rect 130 10531 1580 10542
rect 130 10490 1580 10501
rect 130 10456 138 10490
rect 1572 10456 1580 10490
rect 130 10445 1580 10456
rect 130 10404 1580 10415
rect 130 10370 138 10404
rect 1572 10370 1580 10404
rect 130 10359 1580 10370
rect 130 10318 1580 10329
rect 130 10284 138 10318
rect 1572 10284 1580 10318
rect 130 10273 1580 10284
rect 130 10232 1580 10243
rect 130 10198 138 10232
rect 1572 10198 1580 10232
rect 130 10187 1580 10198
rect 130 10146 1580 10157
rect 130 10112 138 10146
rect 1572 10112 1580 10146
rect 130 10101 1580 10112
rect 130 10060 1580 10071
rect 130 10026 138 10060
rect 1572 10026 1580 10060
rect 130 10015 1580 10026
rect 130 9974 1580 9985
rect 130 9940 138 9974
rect 1572 9940 1580 9974
rect 130 9929 1580 9940
rect 130 9888 1580 9899
rect 130 9854 138 9888
rect 1572 9854 1580 9888
rect 130 9843 1580 9854
rect 130 9802 1580 9813
rect 130 9768 138 9802
rect 1572 9768 1580 9802
rect 130 9757 1580 9768
rect 130 9716 1580 9727
rect 130 9682 138 9716
rect 1572 9682 1580 9716
rect 130 9671 1580 9682
rect 130 9630 1580 9641
rect 130 9596 138 9630
rect 1572 9596 1580 9630
rect 130 9585 1580 9596
rect 130 9544 1580 9555
rect 130 9510 138 9544
rect 1572 9510 1580 9544
rect 130 9499 1580 9510
rect 130 9458 1580 9469
rect 130 9424 138 9458
rect 1572 9424 1580 9458
rect 130 9413 1580 9424
rect 130 9372 1580 9383
rect 130 9338 138 9372
rect 1572 9338 1580 9372
rect 130 9327 1580 9338
rect 130 9286 1580 9297
rect 130 9252 138 9286
rect 1572 9252 1580 9286
rect 130 9241 1580 9252
rect 130 9200 1580 9211
rect 130 9166 138 9200
rect 1572 9166 1580 9200
rect 130 9155 1580 9166
rect 130 9114 1580 9125
rect 130 9080 138 9114
rect 1572 9080 1580 9114
rect 130 9069 1580 9080
rect 130 9028 1580 9039
rect 130 8994 138 9028
rect 1572 8994 1580 9028
rect 130 8983 1580 8994
rect 130 8942 1580 8953
rect 130 8908 138 8942
rect 1572 8908 1580 8942
rect 130 8897 1580 8908
rect 130 8856 1580 8867
rect 130 8822 138 8856
rect 1572 8822 1580 8856
rect 130 8811 1580 8822
rect 130 8770 1580 8781
rect 130 8736 138 8770
rect 1572 8736 1580 8770
rect 130 8725 1580 8736
rect 130 8684 1580 8695
rect 130 8650 138 8684
rect 1572 8650 1580 8684
rect 130 8639 1580 8650
rect 130 8598 1580 8609
rect 130 8564 138 8598
rect 1572 8564 1580 8598
rect 130 8553 1580 8564
rect 130 8512 1580 8523
rect 130 8478 138 8512
rect 1572 8478 1580 8512
rect 130 8467 1580 8478
rect 130 8426 1580 8437
rect 130 8392 138 8426
rect 1572 8392 1580 8426
rect 130 8381 1580 8392
rect 130 8340 1580 8351
rect 130 8306 138 8340
rect 1572 8306 1580 8340
rect 130 8295 1580 8306
rect 130 8254 1580 8265
rect 130 8220 138 8254
rect 1572 8220 1580 8254
rect 130 8209 1580 8220
rect 130 8168 1580 8179
rect 130 8134 138 8168
rect 1572 8134 1580 8168
rect 130 8123 1580 8134
rect 130 8082 1580 8093
rect 130 8048 138 8082
rect 1572 8048 1580 8082
rect 130 8037 1580 8048
rect 130 7996 1580 8007
rect 130 7962 138 7996
rect 1572 7962 1580 7996
rect 130 7951 1580 7962
rect 130 7910 1580 7921
rect 130 7876 138 7910
rect 1572 7876 1580 7910
rect 130 7865 1580 7876
rect 130 7824 1580 7835
rect 130 7790 138 7824
rect 1572 7790 1580 7824
rect 130 7779 1580 7790
rect 130 7738 1580 7749
rect 130 7704 138 7738
rect 1572 7704 1580 7738
rect 130 7693 1580 7704
rect 130 7652 1580 7663
rect 130 7618 138 7652
rect 1572 7618 1580 7652
rect 130 7607 1580 7618
rect 130 7566 1580 7577
rect 130 7532 138 7566
rect 1572 7532 1580 7566
rect 130 7521 1580 7532
rect 130 7480 1580 7491
rect 130 7446 138 7480
rect 1572 7446 1580 7480
rect 130 7435 1580 7446
rect 130 7394 1580 7405
rect 130 7360 138 7394
rect 1572 7360 1580 7394
rect 130 7349 1580 7360
rect 130 7308 1580 7319
rect 130 7274 138 7308
rect 1572 7274 1580 7308
rect 130 7263 1580 7274
rect 130 7222 1580 7233
rect 130 7188 138 7222
rect 1572 7188 1580 7222
rect 130 7177 1580 7188
rect 130 7136 1580 7147
rect 130 7102 138 7136
rect 1572 7102 1580 7136
rect 130 7091 1580 7102
rect 130 7050 1580 7061
rect 130 7016 138 7050
rect 1572 7016 1580 7050
rect 130 7005 1580 7016
rect 130 6964 1580 6975
rect 130 6930 138 6964
rect 1572 6930 1580 6964
rect 130 6919 1580 6930
rect 130 6878 1580 6889
rect 130 6844 138 6878
rect 1572 6844 1580 6878
rect 130 6833 1580 6844
rect 130 6792 1580 6803
rect 130 6758 138 6792
rect 1572 6758 1580 6792
rect 130 6747 1580 6758
rect 130 6706 1580 6717
rect 130 6672 138 6706
rect 1572 6672 1580 6706
rect 130 6661 1580 6672
rect 130 6620 1580 6631
rect 130 6586 138 6620
rect 1572 6586 1580 6620
rect 130 6575 1580 6586
rect 130 6534 1580 6545
rect 130 6500 138 6534
rect 1572 6500 1580 6534
rect 130 6489 1580 6500
rect 130 6448 1580 6459
rect 130 6414 138 6448
rect 1572 6414 1580 6448
rect 130 6403 1580 6414
rect 130 6362 1580 6373
rect 130 6328 138 6362
rect 1572 6328 1580 6362
rect 130 6317 1580 6328
rect 130 6276 1580 6287
rect 130 6242 138 6276
rect 1572 6242 1580 6276
rect 130 6231 1580 6242
rect 130 6190 1580 6201
rect 130 6156 138 6190
rect 1572 6156 1580 6190
rect 130 6145 1580 6156
rect 130 6104 1580 6115
rect 130 6070 138 6104
rect 1572 6070 1580 6104
rect 130 6059 1580 6070
rect 130 6018 1580 6029
rect 130 5984 138 6018
rect 1572 5984 1580 6018
rect 130 5973 1580 5984
rect 130 5932 1580 5943
rect 130 5898 138 5932
rect 1572 5898 1580 5932
rect 130 5887 1580 5898
rect 130 5846 1580 5857
rect 130 5812 138 5846
rect 1572 5812 1580 5846
rect 130 5801 1580 5812
rect 130 5760 1580 5771
rect 130 5726 138 5760
rect 1572 5726 1580 5760
rect 130 5715 1580 5726
rect 130 5674 1580 5685
rect 130 5640 138 5674
rect 1572 5640 1580 5674
rect 130 5629 1580 5640
rect 130 5588 1580 5599
rect 130 5554 138 5588
rect 1572 5554 1580 5588
rect 130 5543 1580 5554
rect 130 5502 1580 5513
rect 130 5468 138 5502
rect 1572 5468 1580 5502
rect 130 5457 1580 5468
rect 130 5416 1580 5427
rect 130 5382 138 5416
rect 1572 5382 1580 5416
rect 130 5371 1580 5382
rect 130 5330 1580 5341
rect 130 5296 138 5330
rect 1572 5296 1580 5330
rect 130 5285 1580 5296
rect 130 5244 1580 5255
rect 130 5210 138 5244
rect 1572 5210 1580 5244
rect 130 5199 1580 5210
rect 130 5158 1580 5169
rect 130 5124 138 5158
rect 1572 5124 1580 5158
rect 130 5113 1580 5124
rect 130 5072 1580 5083
rect 130 5038 138 5072
rect 1572 5038 1580 5072
rect 130 5027 1580 5038
rect 130 4986 1580 4997
rect 130 4952 138 4986
rect 1572 4952 1580 4986
rect 130 4941 1580 4952
rect 130 4900 1580 4911
rect 130 4866 138 4900
rect 1572 4866 1580 4900
rect 130 4855 1580 4866
rect 130 4814 1580 4825
rect 130 4780 138 4814
rect 1572 4780 1580 4814
rect 130 4769 1580 4780
rect 130 4728 1580 4739
rect 130 4694 138 4728
rect 1572 4694 1580 4728
rect 130 4683 1580 4694
rect 130 4642 1580 4653
rect 130 4608 138 4642
rect 1572 4608 1580 4642
rect 130 4597 1580 4608
rect 130 4556 1580 4567
rect 130 4522 138 4556
rect 1572 4522 1580 4556
rect 130 4511 1580 4522
rect 130 4470 1580 4481
rect 130 4436 138 4470
rect 1572 4436 1580 4470
rect 130 4425 1580 4436
rect 130 4384 1580 4395
rect 130 4350 138 4384
rect 1572 4350 1580 4384
rect 130 4339 1580 4350
rect 130 4298 1580 4309
rect 130 4264 138 4298
rect 1572 4264 1580 4298
rect 130 4253 1580 4264
rect 130 4212 1580 4223
rect 130 4178 138 4212
rect 1572 4178 1580 4212
rect 130 4167 1580 4178
rect 130 4126 1580 4137
rect 130 4092 138 4126
rect 1572 4092 1580 4126
rect 130 4081 1580 4092
rect 130 4040 1580 4051
rect 130 4006 138 4040
rect 1572 4006 1580 4040
rect 130 3995 1580 4006
rect 130 3954 1580 3965
rect 130 3920 138 3954
rect 1572 3920 1580 3954
rect 130 3909 1580 3920
rect 130 3868 1580 3879
rect 130 3834 138 3868
rect 1572 3834 1580 3868
rect 130 3823 1580 3834
rect 130 3782 1580 3793
rect 130 3748 138 3782
rect 1572 3748 1580 3782
rect 130 3737 1580 3748
rect 130 3696 1580 3707
rect 130 3662 138 3696
rect 1572 3662 1580 3696
rect 130 3651 1580 3662
rect 130 3610 1580 3621
rect 130 3576 138 3610
rect 1572 3576 1580 3610
rect 130 3565 1580 3576
rect 130 3524 1580 3535
rect 130 3490 138 3524
rect 1572 3490 1580 3524
rect 130 3479 1580 3490
rect 130 3438 1580 3449
rect 130 3404 138 3438
rect 1572 3404 1580 3438
rect 130 3393 1580 3404
rect 130 3352 1580 3363
rect 130 3318 138 3352
rect 1572 3318 1580 3352
rect 130 3307 1580 3318
rect 130 3266 1580 3277
rect 130 3232 138 3266
rect 1572 3232 1580 3266
rect 130 3221 1580 3232
rect 130 3180 1580 3191
rect 130 3146 138 3180
rect 1572 3146 1580 3180
rect 130 3135 1580 3146
rect 130 3094 1580 3105
rect 130 3060 138 3094
rect 1572 3060 1580 3094
rect 130 3049 1580 3060
rect 130 3008 1580 3019
rect 130 2974 138 3008
rect 1572 2974 1580 3008
rect 130 2963 1580 2974
rect 130 2922 1580 2933
rect 130 2888 138 2922
rect 1572 2888 1580 2922
rect 130 2877 1580 2888
rect 130 2836 1580 2847
rect 130 2802 138 2836
rect 1572 2802 1580 2836
rect 130 2791 1580 2802
rect 130 2750 1580 2761
rect 130 2716 138 2750
rect 1572 2716 1580 2750
rect 130 2705 1580 2716
rect 130 2664 1580 2675
rect 130 2630 138 2664
rect 1572 2630 1580 2664
rect 130 2619 1580 2630
rect 130 2578 1580 2589
rect 130 2544 138 2578
rect 1572 2544 1580 2578
rect 130 2533 1580 2544
rect 130 2492 1580 2503
rect 130 2458 138 2492
rect 1572 2458 1580 2492
rect 130 2447 1580 2458
rect 130 2406 1580 2417
rect 130 2372 138 2406
rect 1572 2372 1580 2406
rect 130 2361 1580 2372
rect 130 2320 1580 2331
rect 130 2286 138 2320
rect 1572 2286 1580 2320
rect 130 2275 1580 2286
rect 130 2234 1580 2245
rect 130 2200 138 2234
rect 1572 2200 1580 2234
rect 130 2189 1580 2200
rect 130 2148 1580 2159
rect 130 2114 138 2148
rect 1572 2114 1580 2148
rect 130 2103 1580 2114
rect 130 2062 1580 2073
rect 130 2028 138 2062
rect 1572 2028 1580 2062
rect 130 2017 1580 2028
rect 130 1976 1580 1987
rect 130 1942 138 1976
rect 1572 1942 1580 1976
rect 130 1931 1580 1942
rect 130 1890 1580 1901
rect 130 1856 138 1890
rect 1572 1856 1580 1890
rect 130 1845 1580 1856
rect 130 1804 1580 1815
rect 130 1770 138 1804
rect 1572 1770 1580 1804
rect 130 1759 1580 1770
rect 130 1718 1580 1729
rect 130 1684 138 1718
rect 1572 1684 1580 1718
rect 130 1673 1580 1684
rect 130 1632 1580 1643
rect 130 1598 138 1632
rect 1572 1598 1580 1632
rect 130 1587 1580 1598
rect 130 1546 1580 1557
rect 130 1512 138 1546
rect 1572 1512 1580 1546
rect 130 1501 1580 1512
rect 130 1460 1580 1471
rect 130 1426 138 1460
rect 1572 1426 1580 1460
rect 130 1415 1580 1426
rect 130 1374 1580 1385
rect 130 1340 138 1374
rect 1572 1340 1580 1374
rect 130 1329 1580 1340
rect 130 1288 1580 1299
rect 130 1254 138 1288
rect 1572 1254 1580 1288
rect 130 1243 1580 1254
rect 130 1202 1580 1213
rect 130 1168 138 1202
rect 1572 1168 1580 1202
rect 130 1157 1580 1168
rect 130 1116 1580 1127
rect 130 1082 138 1116
rect 1572 1082 1580 1116
rect 130 1071 1580 1082
rect 130 1030 1580 1041
rect 130 996 138 1030
rect 1572 996 1580 1030
rect 130 985 1580 996
rect 130 944 1580 955
rect 130 910 138 944
rect 1572 910 1580 944
rect 130 899 1580 910
rect 130 858 1580 869
rect 130 824 138 858
rect 1572 824 1580 858
rect 130 813 1580 824
rect 130 772 1580 783
rect 130 738 138 772
rect 1572 738 1580 772
rect 130 727 1580 738
rect 130 686 1580 697
rect 130 652 138 686
rect 1572 652 1580 686
rect 130 641 1580 652
rect 130 600 1580 611
rect 130 566 138 600
rect 1572 566 1580 600
rect 130 555 1580 566
rect 130 514 1580 525
rect 130 480 138 514
rect 1572 480 1580 514
rect 130 469 1580 480
rect 130 428 1580 439
rect 130 394 138 428
rect 1572 394 1580 428
rect 130 383 1580 394
rect 130 342 1580 353
rect 130 308 138 342
rect 1572 308 1580 342
rect 130 297 1580 308
rect 130 256 1580 267
rect 130 222 138 256
rect 1572 222 1580 256
rect 130 211 1580 222
rect 130 170 1580 181
rect 130 136 138 170
rect 1572 136 1580 170
rect 130 124 1580 136
<< pdiffc >>
rect 138 43824 1572 43858
rect 138 43738 1572 43772
rect 138 43652 1572 43686
rect 138 43566 1572 43600
rect 138 43480 1572 43514
rect 138 43394 1572 43428
rect 138 43308 1572 43342
rect 138 43222 1572 43256
rect 138 43136 1572 43170
rect 138 43050 1572 43084
rect 138 42964 1572 42998
rect 138 42878 1572 42912
rect 138 42792 1572 42826
rect 138 42706 1572 42740
rect 138 42620 1572 42654
rect 138 42534 1572 42568
rect 138 42448 1572 42482
rect 138 42362 1572 42396
rect 138 42276 1572 42310
rect 138 42190 1572 42224
rect 138 42104 1572 42138
rect 138 42018 1572 42052
rect 138 41932 1572 41966
rect 138 41846 1572 41880
rect 138 41760 1572 41794
rect 138 41674 1572 41708
rect 138 41588 1572 41622
rect 138 41502 1572 41536
rect 138 41416 1572 41450
rect 138 41330 1572 41364
rect 138 41244 1572 41278
rect 138 41158 1572 41192
rect 138 41072 1572 41106
rect 138 40986 1572 41020
rect 138 40900 1572 40934
rect 138 40814 1572 40848
rect 138 40728 1572 40762
rect 138 40642 1572 40676
rect 138 40556 1572 40590
rect 138 40470 1572 40504
rect 138 40384 1572 40418
rect 138 40298 1572 40332
rect 138 40212 1572 40246
rect 138 40126 1572 40160
rect 138 40040 1572 40074
rect 138 39954 1572 39988
rect 138 39868 1572 39902
rect 138 39782 1572 39816
rect 138 39696 1572 39730
rect 138 39610 1572 39644
rect 138 39524 1572 39558
rect 138 39438 1572 39472
rect 138 39352 1572 39386
rect 138 39266 1572 39300
rect 138 39180 1572 39214
rect 138 39094 1572 39128
rect 138 39008 1572 39042
rect 138 38922 1572 38956
rect 138 38836 1572 38870
rect 138 38750 1572 38784
rect 138 38664 1572 38698
rect 138 38578 1572 38612
rect 138 38492 1572 38526
rect 138 38406 1572 38440
rect 138 38320 1572 38354
rect 138 38234 1572 38268
rect 138 38148 1572 38182
rect 138 38062 1572 38096
rect 138 37976 1572 38010
rect 138 37890 1572 37924
rect 138 37804 1572 37838
rect 138 37718 1572 37752
rect 138 37632 1572 37666
rect 138 37546 1572 37580
rect 138 37460 1572 37494
rect 138 37374 1572 37408
rect 138 37288 1572 37322
rect 138 37202 1572 37236
rect 138 37116 1572 37150
rect 138 37030 1572 37064
rect 138 36944 1572 36978
rect 138 36858 1572 36892
rect 138 36772 1572 36806
rect 138 36686 1572 36720
rect 138 36600 1572 36634
rect 138 36514 1572 36548
rect 138 36428 1572 36462
rect 138 36342 1572 36376
rect 138 36256 1572 36290
rect 138 36170 1572 36204
rect 138 36084 1572 36118
rect 138 35998 1572 36032
rect 138 35912 1572 35946
rect 138 35826 1572 35860
rect 138 35740 1572 35774
rect 138 35654 1572 35688
rect 138 35568 1572 35602
rect 138 35482 1572 35516
rect 138 35396 1572 35430
rect 138 35310 1572 35344
rect 138 35224 1572 35258
rect 138 35138 1572 35172
rect 138 35052 1572 35086
rect 138 34966 1572 35000
rect 138 34880 1572 34914
rect 138 34794 1572 34828
rect 138 34708 1572 34742
rect 138 34622 1572 34656
rect 138 34536 1572 34570
rect 138 34450 1572 34484
rect 138 34364 1572 34398
rect 138 34278 1572 34312
rect 138 34192 1572 34226
rect 138 34106 1572 34140
rect 138 34020 1572 34054
rect 138 33934 1572 33968
rect 138 33848 1572 33882
rect 138 33762 1572 33796
rect 138 33676 1572 33710
rect 138 33590 1572 33624
rect 138 33504 1572 33538
rect 138 33418 1572 33452
rect 138 33332 1572 33366
rect 138 33246 1572 33280
rect 138 33160 1572 33194
rect 138 33074 1572 33108
rect 138 32988 1572 33022
rect 138 32902 1572 32936
rect 138 32816 1572 32850
rect 138 32730 1572 32764
rect 138 32644 1572 32678
rect 138 32558 1572 32592
rect 138 32472 1572 32506
rect 138 32386 1572 32420
rect 138 32300 1572 32334
rect 138 32214 1572 32248
rect 138 32128 1572 32162
rect 138 32042 1572 32076
rect 138 31956 1572 31990
rect 138 31870 1572 31904
rect 138 31784 1572 31818
rect 138 31698 1572 31732
rect 138 31612 1572 31646
rect 138 31526 1572 31560
rect 138 31440 1572 31474
rect 138 31354 1572 31388
rect 138 31268 1572 31302
rect 138 31182 1572 31216
rect 138 31096 1572 31130
rect 138 31010 1572 31044
rect 138 30924 1572 30958
rect 138 30838 1572 30872
rect 138 30752 1572 30786
rect 138 30666 1572 30700
rect 138 30580 1572 30614
rect 138 30494 1572 30528
rect 138 30408 1572 30442
rect 138 30322 1572 30356
rect 138 30236 1572 30270
rect 138 30150 1572 30184
rect 138 30064 1572 30098
rect 138 29978 1572 30012
rect 138 29892 1572 29926
rect 138 29806 1572 29840
rect 138 29720 1572 29754
rect 138 29634 1572 29668
rect 138 29548 1572 29582
rect 138 29462 1572 29496
rect 138 29376 1572 29410
rect 138 29290 1572 29324
rect 138 29204 1572 29238
rect 138 29118 1572 29152
rect 138 29032 1572 29066
rect 138 28946 1572 28980
rect 138 28860 1572 28894
rect 138 28774 1572 28808
rect 138 28688 1572 28722
rect 138 28602 1572 28636
rect 138 28516 1572 28550
rect 138 28430 1572 28464
rect 138 28344 1572 28378
rect 138 28258 1572 28292
rect 138 28172 1572 28206
rect 138 28086 1572 28120
rect 138 28000 1572 28034
rect 138 27914 1572 27948
rect 138 27828 1572 27862
rect 138 27742 1572 27776
rect 138 27656 1572 27690
rect 138 27570 1572 27604
rect 138 27484 1572 27518
rect 138 27398 1572 27432
rect 138 27312 1572 27346
rect 138 27226 1572 27260
rect 138 27140 1572 27174
rect 138 27054 1572 27088
rect 138 26968 1572 27002
rect 138 26882 1572 26916
rect 138 26796 1572 26830
rect 138 26710 1572 26744
rect 138 26624 1572 26658
rect 138 26538 1572 26572
rect 138 26452 1572 26486
rect 138 26366 1572 26400
rect 138 26280 1572 26314
rect 138 26194 1572 26228
rect 138 26108 1572 26142
rect 138 26022 1572 26056
rect 138 25936 1572 25970
rect 138 25850 1572 25884
rect 138 25764 1572 25798
rect 138 25678 1572 25712
rect 138 25592 1572 25626
rect 138 25506 1572 25540
rect 138 25420 1572 25454
rect 138 25334 1572 25368
rect 138 25248 1572 25282
rect 138 25162 1572 25196
rect 138 25076 1572 25110
rect 138 24990 1572 25024
rect 138 24904 1572 24938
rect 138 24818 1572 24852
rect 138 24732 1572 24766
rect 138 24646 1572 24680
rect 138 24560 1572 24594
rect 138 24474 1572 24508
rect 138 24388 1572 24422
rect 138 24302 1572 24336
rect 138 24216 1572 24250
rect 138 24130 1572 24164
rect 138 24044 1572 24078
rect 138 23958 1572 23992
rect 138 23872 1572 23906
rect 138 23786 1572 23820
rect 138 23700 1572 23734
rect 138 23614 1572 23648
rect 138 23528 1572 23562
rect 138 23442 1572 23476
rect 138 23356 1572 23390
rect 138 23270 1572 23304
rect 138 23184 1572 23218
rect 138 23098 1572 23132
rect 138 23012 1572 23046
rect 138 22926 1572 22960
rect 138 22840 1572 22874
rect 138 22754 1572 22788
rect 138 22668 1572 22702
rect 138 22582 1572 22616
rect 138 22496 1572 22530
rect 138 22410 1572 22444
rect 138 22324 1572 22358
rect 138 22238 1572 22272
rect 138 22152 1572 22186
rect 138 22066 1572 22100
rect 138 21980 1572 22014
rect 138 21894 1572 21928
rect 138 21808 1572 21842
rect 138 21722 1572 21756
rect 138 21636 1572 21670
rect 138 21550 1572 21584
rect 138 21464 1572 21498
rect 138 21378 1572 21412
rect 138 21292 1572 21326
rect 138 21206 1572 21240
rect 138 21120 1572 21154
rect 138 21034 1572 21068
rect 138 20948 1572 20982
rect 138 20862 1572 20896
rect 138 20776 1572 20810
rect 138 20690 1572 20724
rect 138 20604 1572 20638
rect 138 20518 1572 20552
rect 138 20432 1572 20466
rect 138 20346 1572 20380
rect 138 20260 1572 20294
rect 138 20174 1572 20208
rect 138 20088 1572 20122
rect 138 20002 1572 20036
rect 138 19916 1572 19950
rect 138 19830 1572 19864
rect 138 19744 1572 19778
rect 138 19658 1572 19692
rect 138 19572 1572 19606
rect 138 19486 1572 19520
rect 138 19400 1572 19434
rect 138 19314 1572 19348
rect 138 19228 1572 19262
rect 138 19142 1572 19176
rect 138 19056 1572 19090
rect 138 18970 1572 19004
rect 138 18884 1572 18918
rect 138 18798 1572 18832
rect 138 18712 1572 18746
rect 138 18626 1572 18660
rect 138 18540 1572 18574
rect 138 18454 1572 18488
rect 138 18368 1572 18402
rect 138 18282 1572 18316
rect 138 18196 1572 18230
rect 138 18110 1572 18144
rect 138 18024 1572 18058
rect 138 17938 1572 17972
rect 138 17852 1572 17886
rect 138 17766 1572 17800
rect 138 17680 1572 17714
rect 138 17594 1572 17628
rect 138 17508 1572 17542
rect 138 17422 1572 17456
rect 138 17336 1572 17370
rect 138 17250 1572 17284
rect 138 17164 1572 17198
rect 138 17078 1572 17112
rect 138 16992 1572 17026
rect 138 16906 1572 16940
rect 138 16820 1572 16854
rect 138 16734 1572 16768
rect 138 16648 1572 16682
rect 138 16562 1572 16596
rect 138 16476 1572 16510
rect 138 16390 1572 16424
rect 138 16304 1572 16338
rect 138 16218 1572 16252
rect 138 16132 1572 16166
rect 138 16046 1572 16080
rect 138 15960 1572 15994
rect 138 15874 1572 15908
rect 138 15788 1572 15822
rect 138 15702 1572 15736
rect 138 15616 1572 15650
rect 138 15530 1572 15564
rect 138 15444 1572 15478
rect 138 15358 1572 15392
rect 138 15272 1572 15306
rect 138 15186 1572 15220
rect 138 15100 1572 15134
rect 138 15014 1572 15048
rect 138 14928 1572 14962
rect 138 14842 1572 14876
rect 138 14756 1572 14790
rect 138 14670 1572 14704
rect 138 14584 1572 14618
rect 138 14498 1572 14532
rect 138 14412 1572 14446
rect 138 14326 1572 14360
rect 138 14240 1572 14274
rect 138 14154 1572 14188
rect 138 14068 1572 14102
rect 138 13982 1572 14016
rect 138 13896 1572 13930
rect 138 13810 1572 13844
rect 138 13724 1572 13758
rect 138 13638 1572 13672
rect 138 13552 1572 13586
rect 138 13466 1572 13500
rect 138 13380 1572 13414
rect 138 13294 1572 13328
rect 138 13208 1572 13242
rect 138 13122 1572 13156
rect 138 13036 1572 13070
rect 138 12950 1572 12984
rect 138 12864 1572 12898
rect 138 12778 1572 12812
rect 138 12692 1572 12726
rect 138 12606 1572 12640
rect 138 12520 1572 12554
rect 138 12434 1572 12468
rect 138 12348 1572 12382
rect 138 12262 1572 12296
rect 138 12176 1572 12210
rect 138 12090 1572 12124
rect 138 12004 1572 12038
rect 138 11918 1572 11952
rect 138 11832 1572 11866
rect 138 11746 1572 11780
rect 138 11660 1572 11694
rect 138 11574 1572 11608
rect 138 11488 1572 11522
rect 138 11402 1572 11436
rect 138 11316 1572 11350
rect 138 11230 1572 11264
rect 138 11144 1572 11178
rect 138 11058 1572 11092
rect 138 10972 1572 11006
rect 138 10886 1572 10920
rect 138 10800 1572 10834
rect 138 10714 1572 10748
rect 138 10628 1572 10662
rect 138 10542 1572 10576
rect 138 10456 1572 10490
rect 138 10370 1572 10404
rect 138 10284 1572 10318
rect 138 10198 1572 10232
rect 138 10112 1572 10146
rect 138 10026 1572 10060
rect 138 9940 1572 9974
rect 138 9854 1572 9888
rect 138 9768 1572 9802
rect 138 9682 1572 9716
rect 138 9596 1572 9630
rect 138 9510 1572 9544
rect 138 9424 1572 9458
rect 138 9338 1572 9372
rect 138 9252 1572 9286
rect 138 9166 1572 9200
rect 138 9080 1572 9114
rect 138 8994 1572 9028
rect 138 8908 1572 8942
rect 138 8822 1572 8856
rect 138 8736 1572 8770
rect 138 8650 1572 8684
rect 138 8564 1572 8598
rect 138 8478 1572 8512
rect 138 8392 1572 8426
rect 138 8306 1572 8340
rect 138 8220 1572 8254
rect 138 8134 1572 8168
rect 138 8048 1572 8082
rect 138 7962 1572 7996
rect 138 7876 1572 7910
rect 138 7790 1572 7824
rect 138 7704 1572 7738
rect 138 7618 1572 7652
rect 138 7532 1572 7566
rect 138 7446 1572 7480
rect 138 7360 1572 7394
rect 138 7274 1572 7308
rect 138 7188 1572 7222
rect 138 7102 1572 7136
rect 138 7016 1572 7050
rect 138 6930 1572 6964
rect 138 6844 1572 6878
rect 138 6758 1572 6792
rect 138 6672 1572 6706
rect 138 6586 1572 6620
rect 138 6500 1572 6534
rect 138 6414 1572 6448
rect 138 6328 1572 6362
rect 138 6242 1572 6276
rect 138 6156 1572 6190
rect 138 6070 1572 6104
rect 138 5984 1572 6018
rect 138 5898 1572 5932
rect 138 5812 1572 5846
rect 138 5726 1572 5760
rect 138 5640 1572 5674
rect 138 5554 1572 5588
rect 138 5468 1572 5502
rect 138 5382 1572 5416
rect 138 5296 1572 5330
rect 138 5210 1572 5244
rect 138 5124 1572 5158
rect 138 5038 1572 5072
rect 138 4952 1572 4986
rect 138 4866 1572 4900
rect 138 4780 1572 4814
rect 138 4694 1572 4728
rect 138 4608 1572 4642
rect 138 4522 1572 4556
rect 138 4436 1572 4470
rect 138 4350 1572 4384
rect 138 4264 1572 4298
rect 138 4178 1572 4212
rect 138 4092 1572 4126
rect 138 4006 1572 4040
rect 138 3920 1572 3954
rect 138 3834 1572 3868
rect 138 3748 1572 3782
rect 138 3662 1572 3696
rect 138 3576 1572 3610
rect 138 3490 1572 3524
rect 138 3404 1572 3438
rect 138 3318 1572 3352
rect 138 3232 1572 3266
rect 138 3146 1572 3180
rect 138 3060 1572 3094
rect 138 2974 1572 3008
rect 138 2888 1572 2922
rect 138 2802 1572 2836
rect 138 2716 1572 2750
rect 138 2630 1572 2664
rect 138 2544 1572 2578
rect 138 2458 1572 2492
rect 138 2372 1572 2406
rect 138 2286 1572 2320
rect 138 2200 1572 2234
rect 138 2114 1572 2148
rect 138 2028 1572 2062
rect 138 1942 1572 1976
rect 138 1856 1572 1890
rect 138 1770 1572 1804
rect 138 1684 1572 1718
rect 138 1598 1572 1632
rect 138 1512 1572 1546
rect 138 1426 1572 1460
rect 138 1340 1572 1374
rect 138 1254 1572 1288
rect 138 1168 1572 1202
rect 138 1082 1572 1116
rect 138 996 1572 1030
rect 138 910 1572 944
rect 138 824 1572 858
rect 138 738 1572 772
rect 138 652 1572 686
rect 138 566 1572 600
rect 138 480 1572 514
rect 138 394 1572 428
rect 138 308 1572 342
rect 138 222 1572 256
rect 138 136 1572 170
<< nsubdiff >>
rect 36 43924 100 43958
rect 1680 43924 1744 43958
rect 36 43894 70 43924
rect 1710 43894 1744 43924
rect 36 70 70 100
rect 1710 70 1744 100
rect 36 36 100 70
rect 1680 36 1744 70
<< nsubdiffcont >>
rect 100 43924 1680 43958
rect 36 100 70 43894
rect 1710 100 1744 43894
rect 100 36 1680 70
<< poly >>
rect 1618 43815 1672 43831
rect 1618 43813 1628 43815
rect 104 43783 130 43813
rect 1580 43783 1628 43813
rect 1618 43727 1628 43783
rect 104 43697 130 43727
rect 1580 43697 1628 43727
rect 1618 43641 1628 43697
rect 104 43611 130 43641
rect 1580 43611 1628 43641
rect 1618 43555 1628 43611
rect 104 43525 130 43555
rect 1580 43525 1628 43555
rect 1618 43469 1628 43525
rect 104 43439 130 43469
rect 1580 43439 1628 43469
rect 1618 43383 1628 43439
rect 104 43353 130 43383
rect 1580 43353 1628 43383
rect 1618 43297 1628 43353
rect 104 43267 130 43297
rect 1580 43267 1628 43297
rect 1618 43211 1628 43267
rect 104 43181 130 43211
rect 1580 43181 1628 43211
rect 1618 43125 1628 43181
rect 104 43095 130 43125
rect 1580 43095 1628 43125
rect 1618 43039 1628 43095
rect 104 43009 130 43039
rect 1580 43009 1628 43039
rect 1618 42953 1628 43009
rect 104 42923 130 42953
rect 1580 42923 1628 42953
rect 1618 42867 1628 42923
rect 104 42837 130 42867
rect 1580 42837 1628 42867
rect 1618 42781 1628 42837
rect 104 42751 130 42781
rect 1580 42751 1628 42781
rect 1618 42695 1628 42751
rect 104 42665 130 42695
rect 1580 42665 1628 42695
rect 1618 42609 1628 42665
rect 104 42579 130 42609
rect 1580 42579 1628 42609
rect 1618 42523 1628 42579
rect 104 42493 130 42523
rect 1580 42493 1628 42523
rect 1618 42437 1628 42493
rect 104 42407 130 42437
rect 1580 42407 1628 42437
rect 1618 42351 1628 42407
rect 104 42321 130 42351
rect 1580 42321 1628 42351
rect 1618 42265 1628 42321
rect 104 42235 130 42265
rect 1580 42235 1628 42265
rect 1618 42179 1628 42235
rect 104 42149 130 42179
rect 1580 42149 1628 42179
rect 1618 42093 1628 42149
rect 104 42063 130 42093
rect 1580 42063 1628 42093
rect 1618 42007 1628 42063
rect 104 41977 130 42007
rect 1580 41977 1628 42007
rect 1618 41921 1628 41977
rect 104 41891 130 41921
rect 1580 41891 1628 41921
rect 1618 41835 1628 41891
rect 104 41805 130 41835
rect 1580 41805 1628 41835
rect 1618 41749 1628 41805
rect 104 41719 130 41749
rect 1580 41719 1628 41749
rect 1618 41663 1628 41719
rect 104 41633 130 41663
rect 1580 41633 1628 41663
rect 1618 41577 1628 41633
rect 104 41547 130 41577
rect 1580 41547 1628 41577
rect 1618 41491 1628 41547
rect 104 41461 130 41491
rect 1580 41461 1628 41491
rect 1618 41405 1628 41461
rect 104 41375 130 41405
rect 1580 41375 1628 41405
rect 1618 41319 1628 41375
rect 104 41289 130 41319
rect 1580 41289 1628 41319
rect 1618 41233 1628 41289
rect 104 41203 130 41233
rect 1580 41203 1628 41233
rect 1618 41147 1628 41203
rect 104 41117 130 41147
rect 1580 41117 1628 41147
rect 1618 41061 1628 41117
rect 104 41031 130 41061
rect 1580 41031 1628 41061
rect 1618 40975 1628 41031
rect 104 40945 130 40975
rect 1580 40945 1628 40975
rect 1618 40889 1628 40945
rect 104 40859 130 40889
rect 1580 40859 1628 40889
rect 1618 40803 1628 40859
rect 104 40773 130 40803
rect 1580 40773 1628 40803
rect 1618 40717 1628 40773
rect 104 40687 130 40717
rect 1580 40687 1628 40717
rect 1618 40631 1628 40687
rect 104 40601 130 40631
rect 1580 40601 1628 40631
rect 1618 40545 1628 40601
rect 104 40515 130 40545
rect 1580 40515 1628 40545
rect 1618 40459 1628 40515
rect 104 40429 130 40459
rect 1580 40429 1628 40459
rect 1618 40373 1628 40429
rect 104 40343 130 40373
rect 1580 40343 1628 40373
rect 1618 40287 1628 40343
rect 104 40257 130 40287
rect 1580 40257 1628 40287
rect 1618 40201 1628 40257
rect 104 40171 130 40201
rect 1580 40171 1628 40201
rect 1618 40115 1628 40171
rect 104 40085 130 40115
rect 1580 40085 1628 40115
rect 1618 40029 1628 40085
rect 104 39999 130 40029
rect 1580 39999 1628 40029
rect 1618 39943 1628 39999
rect 104 39913 130 39943
rect 1580 39913 1628 39943
rect 1618 39857 1628 39913
rect 104 39827 130 39857
rect 1580 39827 1628 39857
rect 1618 39771 1628 39827
rect 104 39741 130 39771
rect 1580 39741 1628 39771
rect 1618 39685 1628 39741
rect 104 39655 130 39685
rect 1580 39655 1628 39685
rect 1618 39599 1628 39655
rect 104 39569 130 39599
rect 1580 39569 1628 39599
rect 1618 39513 1628 39569
rect 104 39483 130 39513
rect 1580 39483 1628 39513
rect 1618 39427 1628 39483
rect 104 39397 130 39427
rect 1580 39397 1628 39427
rect 1618 39341 1628 39397
rect 104 39311 130 39341
rect 1580 39311 1628 39341
rect 1618 39255 1628 39311
rect 104 39225 130 39255
rect 1580 39225 1628 39255
rect 1618 39169 1628 39225
rect 104 39139 130 39169
rect 1580 39139 1628 39169
rect 1618 39083 1628 39139
rect 104 39053 130 39083
rect 1580 39053 1628 39083
rect 1618 38997 1628 39053
rect 104 38967 130 38997
rect 1580 38967 1628 38997
rect 1618 38911 1628 38967
rect 104 38881 130 38911
rect 1580 38881 1628 38911
rect 1618 38825 1628 38881
rect 104 38795 130 38825
rect 1580 38795 1628 38825
rect 1618 38739 1628 38795
rect 104 38709 130 38739
rect 1580 38709 1628 38739
rect 1618 38653 1628 38709
rect 104 38623 130 38653
rect 1580 38623 1628 38653
rect 1618 38567 1628 38623
rect 104 38537 130 38567
rect 1580 38537 1628 38567
rect 1618 38481 1628 38537
rect 104 38451 130 38481
rect 1580 38451 1628 38481
rect 1618 38395 1628 38451
rect 104 38365 130 38395
rect 1580 38365 1628 38395
rect 1618 38309 1628 38365
rect 104 38279 130 38309
rect 1580 38279 1628 38309
rect 1618 38223 1628 38279
rect 104 38193 130 38223
rect 1580 38193 1628 38223
rect 1618 38137 1628 38193
rect 104 38107 130 38137
rect 1580 38107 1628 38137
rect 1618 38051 1628 38107
rect 104 38021 130 38051
rect 1580 38021 1628 38051
rect 1618 37965 1628 38021
rect 104 37935 130 37965
rect 1580 37935 1628 37965
rect 1618 37879 1628 37935
rect 104 37849 130 37879
rect 1580 37849 1628 37879
rect 1618 37793 1628 37849
rect 104 37763 130 37793
rect 1580 37763 1628 37793
rect 1618 37707 1628 37763
rect 104 37677 130 37707
rect 1580 37677 1628 37707
rect 1618 37621 1628 37677
rect 104 37591 130 37621
rect 1580 37591 1628 37621
rect 1618 37535 1628 37591
rect 104 37505 130 37535
rect 1580 37505 1628 37535
rect 1618 37449 1628 37505
rect 104 37419 130 37449
rect 1580 37419 1628 37449
rect 1618 37363 1628 37419
rect 104 37333 130 37363
rect 1580 37333 1628 37363
rect 1618 37277 1628 37333
rect 104 37247 130 37277
rect 1580 37247 1628 37277
rect 1618 37191 1628 37247
rect 104 37161 130 37191
rect 1580 37161 1628 37191
rect 1618 37105 1628 37161
rect 104 37075 130 37105
rect 1580 37075 1628 37105
rect 1618 37019 1628 37075
rect 104 36989 130 37019
rect 1580 36989 1628 37019
rect 1618 36933 1628 36989
rect 104 36903 130 36933
rect 1580 36903 1628 36933
rect 1618 36847 1628 36903
rect 104 36817 130 36847
rect 1580 36817 1628 36847
rect 1618 36761 1628 36817
rect 104 36731 130 36761
rect 1580 36731 1628 36761
rect 1618 36675 1628 36731
rect 104 36645 130 36675
rect 1580 36645 1628 36675
rect 1618 36589 1628 36645
rect 104 36559 130 36589
rect 1580 36559 1628 36589
rect 1618 36503 1628 36559
rect 104 36473 130 36503
rect 1580 36473 1628 36503
rect 1618 36417 1628 36473
rect 104 36387 130 36417
rect 1580 36387 1628 36417
rect 1618 36331 1628 36387
rect 104 36301 130 36331
rect 1580 36301 1628 36331
rect 1618 36245 1628 36301
rect 104 36215 130 36245
rect 1580 36215 1628 36245
rect 1618 36159 1628 36215
rect 104 36129 130 36159
rect 1580 36129 1628 36159
rect 1618 36073 1628 36129
rect 104 36043 130 36073
rect 1580 36043 1628 36073
rect 1618 35987 1628 36043
rect 104 35957 130 35987
rect 1580 35957 1628 35987
rect 1618 35901 1628 35957
rect 104 35871 130 35901
rect 1580 35871 1628 35901
rect 1618 35815 1628 35871
rect 104 35785 130 35815
rect 1580 35785 1628 35815
rect 1618 35729 1628 35785
rect 104 35699 130 35729
rect 1580 35699 1628 35729
rect 1618 35643 1628 35699
rect 104 35613 130 35643
rect 1580 35613 1628 35643
rect 1618 35557 1628 35613
rect 104 35527 130 35557
rect 1580 35527 1628 35557
rect 1618 35471 1628 35527
rect 104 35441 130 35471
rect 1580 35441 1628 35471
rect 1618 35385 1628 35441
rect 104 35355 130 35385
rect 1580 35355 1628 35385
rect 1618 35299 1628 35355
rect 104 35269 130 35299
rect 1580 35269 1628 35299
rect 1618 35213 1628 35269
rect 104 35183 130 35213
rect 1580 35183 1628 35213
rect 1618 35127 1628 35183
rect 104 35097 130 35127
rect 1580 35097 1628 35127
rect 1618 35041 1628 35097
rect 104 35011 130 35041
rect 1580 35011 1628 35041
rect 1618 34955 1628 35011
rect 104 34925 130 34955
rect 1580 34925 1628 34955
rect 1618 34869 1628 34925
rect 104 34839 130 34869
rect 1580 34839 1628 34869
rect 1618 34783 1628 34839
rect 104 34753 130 34783
rect 1580 34753 1628 34783
rect 1618 34697 1628 34753
rect 104 34667 130 34697
rect 1580 34667 1628 34697
rect 1618 34611 1628 34667
rect 104 34581 130 34611
rect 1580 34581 1628 34611
rect 1618 34525 1628 34581
rect 104 34495 130 34525
rect 1580 34495 1628 34525
rect 1618 34439 1628 34495
rect 104 34409 130 34439
rect 1580 34409 1628 34439
rect 1618 34353 1628 34409
rect 104 34323 130 34353
rect 1580 34323 1628 34353
rect 1618 34267 1628 34323
rect 104 34237 130 34267
rect 1580 34237 1628 34267
rect 1618 34181 1628 34237
rect 104 34151 130 34181
rect 1580 34151 1628 34181
rect 1618 34095 1628 34151
rect 104 34065 130 34095
rect 1580 34065 1628 34095
rect 1618 34009 1628 34065
rect 104 33979 130 34009
rect 1580 33979 1628 34009
rect 1618 33923 1628 33979
rect 104 33893 130 33923
rect 1580 33893 1628 33923
rect 1618 33837 1628 33893
rect 104 33807 130 33837
rect 1580 33807 1628 33837
rect 1618 33751 1628 33807
rect 104 33721 130 33751
rect 1580 33721 1628 33751
rect 1618 33665 1628 33721
rect 104 33635 130 33665
rect 1580 33635 1628 33665
rect 1618 33579 1628 33635
rect 104 33549 130 33579
rect 1580 33549 1628 33579
rect 1618 33493 1628 33549
rect 104 33463 130 33493
rect 1580 33463 1628 33493
rect 1618 33407 1628 33463
rect 104 33377 130 33407
rect 1580 33377 1628 33407
rect 1618 33321 1628 33377
rect 104 33291 130 33321
rect 1580 33291 1628 33321
rect 1618 33235 1628 33291
rect 104 33205 130 33235
rect 1580 33205 1628 33235
rect 1618 33149 1628 33205
rect 104 33119 130 33149
rect 1580 33119 1628 33149
rect 1618 33063 1628 33119
rect 104 33033 130 33063
rect 1580 33033 1628 33063
rect 1618 32977 1628 33033
rect 104 32947 130 32977
rect 1580 32947 1628 32977
rect 1618 32891 1628 32947
rect 104 32861 130 32891
rect 1580 32861 1628 32891
rect 1618 32805 1628 32861
rect 104 32775 130 32805
rect 1580 32775 1628 32805
rect 1618 32719 1628 32775
rect 104 32689 130 32719
rect 1580 32689 1628 32719
rect 1618 32633 1628 32689
rect 104 32603 130 32633
rect 1580 32603 1628 32633
rect 1618 32547 1628 32603
rect 104 32517 130 32547
rect 1580 32517 1628 32547
rect 1618 32461 1628 32517
rect 104 32431 130 32461
rect 1580 32431 1628 32461
rect 1618 32375 1628 32431
rect 104 32345 130 32375
rect 1580 32345 1628 32375
rect 1618 32289 1628 32345
rect 104 32259 130 32289
rect 1580 32259 1628 32289
rect 1618 32203 1628 32259
rect 104 32173 130 32203
rect 1580 32173 1628 32203
rect 1618 32117 1628 32173
rect 104 32087 130 32117
rect 1580 32087 1628 32117
rect 1618 32031 1628 32087
rect 104 32001 130 32031
rect 1580 32001 1628 32031
rect 1618 31945 1628 32001
rect 104 31915 130 31945
rect 1580 31915 1628 31945
rect 1618 31859 1628 31915
rect 104 31829 130 31859
rect 1580 31829 1628 31859
rect 1618 31773 1628 31829
rect 104 31743 130 31773
rect 1580 31743 1628 31773
rect 1618 31687 1628 31743
rect 104 31657 130 31687
rect 1580 31657 1628 31687
rect 1618 31601 1628 31657
rect 104 31571 130 31601
rect 1580 31571 1628 31601
rect 1618 31515 1628 31571
rect 104 31485 130 31515
rect 1580 31485 1628 31515
rect 1618 31429 1628 31485
rect 104 31399 130 31429
rect 1580 31399 1628 31429
rect 1618 31343 1628 31399
rect 104 31313 130 31343
rect 1580 31313 1628 31343
rect 1618 31257 1628 31313
rect 104 31227 130 31257
rect 1580 31227 1628 31257
rect 1618 31171 1628 31227
rect 104 31141 130 31171
rect 1580 31141 1628 31171
rect 1618 31085 1628 31141
rect 104 31055 130 31085
rect 1580 31055 1628 31085
rect 1618 30999 1628 31055
rect 104 30969 130 30999
rect 1580 30969 1628 30999
rect 1618 30913 1628 30969
rect 104 30883 130 30913
rect 1580 30883 1628 30913
rect 1618 30827 1628 30883
rect 104 30797 130 30827
rect 1580 30797 1628 30827
rect 1618 30741 1628 30797
rect 104 30711 130 30741
rect 1580 30711 1628 30741
rect 1618 30655 1628 30711
rect 104 30625 130 30655
rect 1580 30625 1628 30655
rect 1618 30569 1628 30625
rect 104 30539 130 30569
rect 1580 30539 1628 30569
rect 1618 30483 1628 30539
rect 104 30453 130 30483
rect 1580 30453 1628 30483
rect 1618 30397 1628 30453
rect 104 30367 130 30397
rect 1580 30367 1628 30397
rect 1618 30311 1628 30367
rect 104 30281 130 30311
rect 1580 30281 1628 30311
rect 1618 30225 1628 30281
rect 104 30195 130 30225
rect 1580 30195 1628 30225
rect 1618 30139 1628 30195
rect 104 30109 130 30139
rect 1580 30109 1628 30139
rect 1618 30053 1628 30109
rect 104 30023 130 30053
rect 1580 30023 1628 30053
rect 1618 29967 1628 30023
rect 104 29937 130 29967
rect 1580 29937 1628 29967
rect 1618 29881 1628 29937
rect 104 29851 130 29881
rect 1580 29851 1628 29881
rect 1618 29795 1628 29851
rect 104 29765 130 29795
rect 1580 29765 1628 29795
rect 1618 29709 1628 29765
rect 104 29679 130 29709
rect 1580 29679 1628 29709
rect 1618 29623 1628 29679
rect 104 29593 130 29623
rect 1580 29593 1628 29623
rect 1618 29537 1628 29593
rect 104 29507 130 29537
rect 1580 29507 1628 29537
rect 1618 29451 1628 29507
rect 104 29421 130 29451
rect 1580 29421 1628 29451
rect 1618 29365 1628 29421
rect 104 29335 130 29365
rect 1580 29335 1628 29365
rect 1618 29279 1628 29335
rect 104 29249 130 29279
rect 1580 29249 1628 29279
rect 1618 29193 1628 29249
rect 104 29163 130 29193
rect 1580 29163 1628 29193
rect 1618 29107 1628 29163
rect 104 29077 130 29107
rect 1580 29077 1628 29107
rect 1618 29021 1628 29077
rect 104 28991 130 29021
rect 1580 28991 1628 29021
rect 1618 28935 1628 28991
rect 104 28905 130 28935
rect 1580 28905 1628 28935
rect 1618 28849 1628 28905
rect 104 28819 130 28849
rect 1580 28819 1628 28849
rect 1618 28763 1628 28819
rect 104 28733 130 28763
rect 1580 28733 1628 28763
rect 1618 28677 1628 28733
rect 104 28647 130 28677
rect 1580 28647 1628 28677
rect 1618 28591 1628 28647
rect 104 28561 130 28591
rect 1580 28561 1628 28591
rect 1618 28505 1628 28561
rect 104 28475 130 28505
rect 1580 28475 1628 28505
rect 1618 28419 1628 28475
rect 104 28389 130 28419
rect 1580 28389 1628 28419
rect 1618 28333 1628 28389
rect 104 28303 130 28333
rect 1580 28303 1628 28333
rect 1618 28247 1628 28303
rect 104 28217 130 28247
rect 1580 28217 1628 28247
rect 1618 28161 1628 28217
rect 104 28131 130 28161
rect 1580 28131 1628 28161
rect 1618 28075 1628 28131
rect 104 28045 130 28075
rect 1580 28045 1628 28075
rect 1618 27989 1628 28045
rect 104 27959 130 27989
rect 1580 27959 1628 27989
rect 1618 27903 1628 27959
rect 104 27873 130 27903
rect 1580 27873 1628 27903
rect 1618 27817 1628 27873
rect 104 27787 130 27817
rect 1580 27787 1628 27817
rect 1618 27731 1628 27787
rect 104 27701 130 27731
rect 1580 27701 1628 27731
rect 1618 27645 1628 27701
rect 104 27615 130 27645
rect 1580 27615 1628 27645
rect 1618 27559 1628 27615
rect 104 27529 130 27559
rect 1580 27529 1628 27559
rect 1618 27473 1628 27529
rect 104 27443 130 27473
rect 1580 27443 1628 27473
rect 1618 27387 1628 27443
rect 104 27357 130 27387
rect 1580 27357 1628 27387
rect 1618 27301 1628 27357
rect 104 27271 130 27301
rect 1580 27271 1628 27301
rect 1618 27215 1628 27271
rect 104 27185 130 27215
rect 1580 27185 1628 27215
rect 1618 27129 1628 27185
rect 104 27099 130 27129
rect 1580 27099 1628 27129
rect 1618 27043 1628 27099
rect 104 27013 130 27043
rect 1580 27013 1628 27043
rect 1618 26957 1628 27013
rect 104 26927 130 26957
rect 1580 26927 1628 26957
rect 1618 26871 1628 26927
rect 104 26841 130 26871
rect 1580 26841 1628 26871
rect 1618 26785 1628 26841
rect 104 26755 130 26785
rect 1580 26755 1628 26785
rect 1618 26699 1628 26755
rect 104 26669 130 26699
rect 1580 26669 1628 26699
rect 1618 26613 1628 26669
rect 104 26583 130 26613
rect 1580 26583 1628 26613
rect 1618 26527 1628 26583
rect 104 26497 130 26527
rect 1580 26497 1628 26527
rect 1618 26441 1628 26497
rect 104 26411 130 26441
rect 1580 26411 1628 26441
rect 1618 26355 1628 26411
rect 104 26325 130 26355
rect 1580 26325 1628 26355
rect 1618 26269 1628 26325
rect 104 26239 130 26269
rect 1580 26239 1628 26269
rect 1618 26183 1628 26239
rect 104 26153 130 26183
rect 1580 26153 1628 26183
rect 1618 26097 1628 26153
rect 104 26067 130 26097
rect 1580 26067 1628 26097
rect 1618 26011 1628 26067
rect 104 25981 130 26011
rect 1580 25981 1628 26011
rect 1618 25925 1628 25981
rect 104 25895 130 25925
rect 1580 25895 1628 25925
rect 1618 25839 1628 25895
rect 104 25809 130 25839
rect 1580 25809 1628 25839
rect 1618 25753 1628 25809
rect 104 25723 130 25753
rect 1580 25723 1628 25753
rect 1618 25667 1628 25723
rect 104 25637 130 25667
rect 1580 25637 1628 25667
rect 1618 25581 1628 25637
rect 104 25551 130 25581
rect 1580 25551 1628 25581
rect 1618 25495 1628 25551
rect 104 25465 130 25495
rect 1580 25465 1628 25495
rect 1618 25409 1628 25465
rect 104 25379 130 25409
rect 1580 25379 1628 25409
rect 1618 25323 1628 25379
rect 104 25293 130 25323
rect 1580 25293 1628 25323
rect 1618 25237 1628 25293
rect 104 25207 130 25237
rect 1580 25207 1628 25237
rect 1618 25151 1628 25207
rect 104 25121 130 25151
rect 1580 25121 1628 25151
rect 1618 25065 1628 25121
rect 104 25035 130 25065
rect 1580 25035 1628 25065
rect 1618 24979 1628 25035
rect 104 24949 130 24979
rect 1580 24949 1628 24979
rect 1618 24893 1628 24949
rect 104 24863 130 24893
rect 1580 24863 1628 24893
rect 1618 24807 1628 24863
rect 104 24777 130 24807
rect 1580 24777 1628 24807
rect 1618 24721 1628 24777
rect 104 24691 130 24721
rect 1580 24691 1628 24721
rect 1618 24635 1628 24691
rect 104 24605 130 24635
rect 1580 24605 1628 24635
rect 1618 24549 1628 24605
rect 104 24519 130 24549
rect 1580 24519 1628 24549
rect 1618 24463 1628 24519
rect 104 24433 130 24463
rect 1580 24433 1628 24463
rect 1618 24377 1628 24433
rect 104 24347 130 24377
rect 1580 24347 1628 24377
rect 1618 24291 1628 24347
rect 104 24261 130 24291
rect 1580 24261 1628 24291
rect 1618 24205 1628 24261
rect 104 24175 130 24205
rect 1580 24175 1628 24205
rect 1618 24119 1628 24175
rect 104 24089 130 24119
rect 1580 24089 1628 24119
rect 1618 24033 1628 24089
rect 104 24003 130 24033
rect 1580 24003 1628 24033
rect 1618 23947 1628 24003
rect 104 23917 130 23947
rect 1580 23917 1628 23947
rect 1618 23861 1628 23917
rect 104 23831 130 23861
rect 1580 23831 1628 23861
rect 1618 23775 1628 23831
rect 104 23745 130 23775
rect 1580 23745 1628 23775
rect 1618 23689 1628 23745
rect 104 23659 130 23689
rect 1580 23659 1628 23689
rect 1618 23603 1628 23659
rect 104 23573 130 23603
rect 1580 23573 1628 23603
rect 1618 23517 1628 23573
rect 104 23487 130 23517
rect 1580 23487 1628 23517
rect 1618 23431 1628 23487
rect 104 23401 130 23431
rect 1580 23401 1628 23431
rect 1618 23345 1628 23401
rect 104 23315 130 23345
rect 1580 23315 1628 23345
rect 1618 23259 1628 23315
rect 104 23229 130 23259
rect 1580 23229 1628 23259
rect 1618 23173 1628 23229
rect 104 23143 130 23173
rect 1580 23143 1628 23173
rect 1618 23087 1628 23143
rect 104 23057 130 23087
rect 1580 23057 1628 23087
rect 1618 23001 1628 23057
rect 104 22971 130 23001
rect 1580 22971 1628 23001
rect 1618 22915 1628 22971
rect 104 22885 130 22915
rect 1580 22885 1628 22915
rect 1618 22829 1628 22885
rect 104 22799 130 22829
rect 1580 22799 1628 22829
rect 1618 22743 1628 22799
rect 104 22713 130 22743
rect 1580 22713 1628 22743
rect 1618 22657 1628 22713
rect 104 22627 130 22657
rect 1580 22627 1628 22657
rect 1618 22571 1628 22627
rect 104 22541 130 22571
rect 1580 22541 1628 22571
rect 1618 22485 1628 22541
rect 104 22455 130 22485
rect 1580 22455 1628 22485
rect 1618 22399 1628 22455
rect 104 22369 130 22399
rect 1580 22369 1628 22399
rect 1618 22313 1628 22369
rect 104 22283 130 22313
rect 1580 22283 1628 22313
rect 1618 22227 1628 22283
rect 104 22197 130 22227
rect 1580 22197 1628 22227
rect 1618 22141 1628 22197
rect 104 22111 130 22141
rect 1580 22111 1628 22141
rect 1618 22055 1628 22111
rect 104 22025 130 22055
rect 1580 22025 1628 22055
rect 1618 21969 1628 22025
rect 104 21939 130 21969
rect 1580 21939 1628 21969
rect 1618 21883 1628 21939
rect 104 21853 130 21883
rect 1580 21853 1628 21883
rect 1618 21797 1628 21853
rect 104 21767 130 21797
rect 1580 21767 1628 21797
rect 1618 21711 1628 21767
rect 104 21681 130 21711
rect 1580 21681 1628 21711
rect 1618 21625 1628 21681
rect 104 21595 130 21625
rect 1580 21595 1628 21625
rect 1618 21539 1628 21595
rect 104 21509 130 21539
rect 1580 21509 1628 21539
rect 1618 21453 1628 21509
rect 104 21423 130 21453
rect 1580 21423 1628 21453
rect 1618 21367 1628 21423
rect 104 21337 130 21367
rect 1580 21337 1628 21367
rect 1618 21281 1628 21337
rect 104 21251 130 21281
rect 1580 21251 1628 21281
rect 1618 21195 1628 21251
rect 104 21165 130 21195
rect 1580 21165 1628 21195
rect 1618 21109 1628 21165
rect 104 21079 130 21109
rect 1580 21079 1628 21109
rect 1618 21023 1628 21079
rect 104 20993 130 21023
rect 1580 20993 1628 21023
rect 1618 20937 1628 20993
rect 104 20907 130 20937
rect 1580 20907 1628 20937
rect 1618 20851 1628 20907
rect 104 20821 130 20851
rect 1580 20821 1628 20851
rect 1618 20765 1628 20821
rect 104 20735 130 20765
rect 1580 20735 1628 20765
rect 1618 20679 1628 20735
rect 104 20649 130 20679
rect 1580 20649 1628 20679
rect 1618 20593 1628 20649
rect 104 20563 130 20593
rect 1580 20563 1628 20593
rect 1618 20507 1628 20563
rect 104 20477 130 20507
rect 1580 20477 1628 20507
rect 1618 20421 1628 20477
rect 104 20391 130 20421
rect 1580 20391 1628 20421
rect 1618 20335 1628 20391
rect 104 20305 130 20335
rect 1580 20305 1628 20335
rect 1618 20249 1628 20305
rect 104 20219 130 20249
rect 1580 20219 1628 20249
rect 1618 20163 1628 20219
rect 104 20133 130 20163
rect 1580 20133 1628 20163
rect 1618 20077 1628 20133
rect 104 20047 130 20077
rect 1580 20047 1628 20077
rect 1618 19991 1628 20047
rect 104 19961 130 19991
rect 1580 19961 1628 19991
rect 1618 19905 1628 19961
rect 104 19875 130 19905
rect 1580 19875 1628 19905
rect 1618 19819 1628 19875
rect 104 19789 130 19819
rect 1580 19789 1628 19819
rect 1618 19733 1628 19789
rect 104 19703 130 19733
rect 1580 19703 1628 19733
rect 1618 19647 1628 19703
rect 104 19617 130 19647
rect 1580 19617 1628 19647
rect 1618 19561 1628 19617
rect 104 19531 130 19561
rect 1580 19531 1628 19561
rect 1618 19475 1628 19531
rect 104 19445 130 19475
rect 1580 19445 1628 19475
rect 1618 19389 1628 19445
rect 104 19359 130 19389
rect 1580 19359 1628 19389
rect 1618 19303 1628 19359
rect 104 19273 130 19303
rect 1580 19273 1628 19303
rect 1618 19217 1628 19273
rect 104 19187 130 19217
rect 1580 19187 1628 19217
rect 1618 19131 1628 19187
rect 104 19101 130 19131
rect 1580 19101 1628 19131
rect 1618 19045 1628 19101
rect 104 19015 130 19045
rect 1580 19015 1628 19045
rect 1618 18959 1628 19015
rect 104 18929 130 18959
rect 1580 18929 1628 18959
rect 1618 18873 1628 18929
rect 104 18843 130 18873
rect 1580 18843 1628 18873
rect 1618 18787 1628 18843
rect 104 18757 130 18787
rect 1580 18757 1628 18787
rect 1618 18701 1628 18757
rect 104 18671 130 18701
rect 1580 18671 1628 18701
rect 1618 18615 1628 18671
rect 104 18585 130 18615
rect 1580 18585 1628 18615
rect 1618 18529 1628 18585
rect 104 18499 130 18529
rect 1580 18499 1628 18529
rect 1618 18443 1628 18499
rect 104 18413 130 18443
rect 1580 18413 1628 18443
rect 1618 18357 1628 18413
rect 104 18327 130 18357
rect 1580 18327 1628 18357
rect 1618 18271 1628 18327
rect 104 18241 130 18271
rect 1580 18241 1628 18271
rect 1618 18185 1628 18241
rect 104 18155 130 18185
rect 1580 18155 1628 18185
rect 1618 18099 1628 18155
rect 104 18069 130 18099
rect 1580 18069 1628 18099
rect 1618 18013 1628 18069
rect 104 17983 130 18013
rect 1580 17983 1628 18013
rect 1618 17927 1628 17983
rect 104 17897 130 17927
rect 1580 17897 1628 17927
rect 1618 17841 1628 17897
rect 104 17811 130 17841
rect 1580 17811 1628 17841
rect 1618 17755 1628 17811
rect 104 17725 130 17755
rect 1580 17725 1628 17755
rect 1618 17669 1628 17725
rect 104 17639 130 17669
rect 1580 17639 1628 17669
rect 1618 17583 1628 17639
rect 104 17553 130 17583
rect 1580 17553 1628 17583
rect 1618 17497 1628 17553
rect 104 17467 130 17497
rect 1580 17467 1628 17497
rect 1618 17411 1628 17467
rect 104 17381 130 17411
rect 1580 17381 1628 17411
rect 1618 17325 1628 17381
rect 104 17295 130 17325
rect 1580 17295 1628 17325
rect 1618 17239 1628 17295
rect 104 17209 130 17239
rect 1580 17209 1628 17239
rect 1618 17153 1628 17209
rect 104 17123 130 17153
rect 1580 17123 1628 17153
rect 1618 17067 1628 17123
rect 104 17037 130 17067
rect 1580 17037 1628 17067
rect 1618 16981 1628 17037
rect 104 16951 130 16981
rect 1580 16951 1628 16981
rect 1618 16895 1628 16951
rect 104 16865 130 16895
rect 1580 16865 1628 16895
rect 1618 16809 1628 16865
rect 104 16779 130 16809
rect 1580 16779 1628 16809
rect 1618 16723 1628 16779
rect 104 16693 130 16723
rect 1580 16693 1628 16723
rect 1618 16637 1628 16693
rect 104 16607 130 16637
rect 1580 16607 1628 16637
rect 1618 16551 1628 16607
rect 104 16521 130 16551
rect 1580 16521 1628 16551
rect 1618 16465 1628 16521
rect 104 16435 130 16465
rect 1580 16435 1628 16465
rect 1618 16379 1628 16435
rect 104 16349 130 16379
rect 1580 16349 1628 16379
rect 1618 16293 1628 16349
rect 104 16263 130 16293
rect 1580 16263 1628 16293
rect 1618 16207 1628 16263
rect 104 16177 130 16207
rect 1580 16177 1628 16207
rect 1618 16121 1628 16177
rect 104 16091 130 16121
rect 1580 16091 1628 16121
rect 1618 16035 1628 16091
rect 104 16005 130 16035
rect 1580 16005 1628 16035
rect 1618 15949 1628 16005
rect 104 15919 130 15949
rect 1580 15919 1628 15949
rect 1618 15863 1628 15919
rect 104 15833 130 15863
rect 1580 15833 1628 15863
rect 1618 15777 1628 15833
rect 104 15747 130 15777
rect 1580 15747 1628 15777
rect 1618 15691 1628 15747
rect 104 15661 130 15691
rect 1580 15661 1628 15691
rect 1618 15605 1628 15661
rect 104 15575 130 15605
rect 1580 15575 1628 15605
rect 1618 15519 1628 15575
rect 104 15489 130 15519
rect 1580 15489 1628 15519
rect 1618 15433 1628 15489
rect 104 15403 130 15433
rect 1580 15403 1628 15433
rect 1618 15347 1628 15403
rect 104 15317 130 15347
rect 1580 15317 1628 15347
rect 1618 15261 1628 15317
rect 104 15231 130 15261
rect 1580 15231 1628 15261
rect 1618 15175 1628 15231
rect 104 15145 130 15175
rect 1580 15145 1628 15175
rect 1618 15089 1628 15145
rect 104 15059 130 15089
rect 1580 15059 1628 15089
rect 1618 15003 1628 15059
rect 104 14973 130 15003
rect 1580 14973 1628 15003
rect 1618 14917 1628 14973
rect 104 14887 130 14917
rect 1580 14887 1628 14917
rect 1618 14831 1628 14887
rect 104 14801 130 14831
rect 1580 14801 1628 14831
rect 1618 14745 1628 14801
rect 104 14715 130 14745
rect 1580 14715 1628 14745
rect 1618 14659 1628 14715
rect 104 14629 130 14659
rect 1580 14629 1628 14659
rect 1618 14573 1628 14629
rect 104 14543 130 14573
rect 1580 14543 1628 14573
rect 1618 14487 1628 14543
rect 104 14457 130 14487
rect 1580 14457 1628 14487
rect 1618 14401 1628 14457
rect 104 14371 130 14401
rect 1580 14371 1628 14401
rect 1618 14315 1628 14371
rect 104 14285 130 14315
rect 1580 14285 1628 14315
rect 1618 14229 1628 14285
rect 104 14199 130 14229
rect 1580 14199 1628 14229
rect 1618 14143 1628 14199
rect 104 14113 130 14143
rect 1580 14113 1628 14143
rect 1618 14057 1628 14113
rect 104 14027 130 14057
rect 1580 14027 1628 14057
rect 1618 13971 1628 14027
rect 104 13941 130 13971
rect 1580 13941 1628 13971
rect 1618 13885 1628 13941
rect 104 13855 130 13885
rect 1580 13855 1628 13885
rect 1618 13799 1628 13855
rect 104 13769 130 13799
rect 1580 13769 1628 13799
rect 1618 13713 1628 13769
rect 104 13683 130 13713
rect 1580 13683 1628 13713
rect 1618 13627 1628 13683
rect 104 13597 130 13627
rect 1580 13597 1628 13627
rect 1618 13541 1628 13597
rect 104 13511 130 13541
rect 1580 13511 1628 13541
rect 1618 13455 1628 13511
rect 104 13425 130 13455
rect 1580 13425 1628 13455
rect 1618 13369 1628 13425
rect 104 13339 130 13369
rect 1580 13339 1628 13369
rect 1618 13283 1628 13339
rect 104 13253 130 13283
rect 1580 13253 1628 13283
rect 1618 13197 1628 13253
rect 104 13167 130 13197
rect 1580 13167 1628 13197
rect 1618 13111 1628 13167
rect 104 13081 130 13111
rect 1580 13081 1628 13111
rect 1618 13025 1628 13081
rect 104 12995 130 13025
rect 1580 12995 1628 13025
rect 1618 12939 1628 12995
rect 104 12909 130 12939
rect 1580 12909 1628 12939
rect 1618 12853 1628 12909
rect 104 12823 130 12853
rect 1580 12823 1628 12853
rect 1618 12767 1628 12823
rect 104 12737 130 12767
rect 1580 12737 1628 12767
rect 1618 12681 1628 12737
rect 104 12651 130 12681
rect 1580 12651 1628 12681
rect 1618 12595 1628 12651
rect 104 12565 130 12595
rect 1580 12565 1628 12595
rect 1618 12509 1628 12565
rect 104 12479 130 12509
rect 1580 12479 1628 12509
rect 1618 12423 1628 12479
rect 104 12393 130 12423
rect 1580 12393 1628 12423
rect 1618 12337 1628 12393
rect 104 12307 130 12337
rect 1580 12307 1628 12337
rect 1618 12251 1628 12307
rect 104 12221 130 12251
rect 1580 12221 1628 12251
rect 1618 12165 1628 12221
rect 104 12135 130 12165
rect 1580 12135 1628 12165
rect 1618 12079 1628 12135
rect 104 12049 130 12079
rect 1580 12049 1628 12079
rect 1618 11993 1628 12049
rect 104 11963 130 11993
rect 1580 11963 1628 11993
rect 1618 11907 1628 11963
rect 104 11877 130 11907
rect 1580 11877 1628 11907
rect 1618 11821 1628 11877
rect 104 11791 130 11821
rect 1580 11791 1628 11821
rect 1618 11735 1628 11791
rect 104 11705 130 11735
rect 1580 11705 1628 11735
rect 1618 11649 1628 11705
rect 104 11619 130 11649
rect 1580 11619 1628 11649
rect 1618 11563 1628 11619
rect 104 11533 130 11563
rect 1580 11533 1628 11563
rect 1618 11477 1628 11533
rect 104 11447 130 11477
rect 1580 11447 1628 11477
rect 1618 11391 1628 11447
rect 104 11361 130 11391
rect 1580 11361 1628 11391
rect 1618 11305 1628 11361
rect 104 11275 130 11305
rect 1580 11275 1628 11305
rect 1618 11219 1628 11275
rect 104 11189 130 11219
rect 1580 11189 1628 11219
rect 1618 11133 1628 11189
rect 104 11103 130 11133
rect 1580 11103 1628 11133
rect 1618 11047 1628 11103
rect 104 11017 130 11047
rect 1580 11017 1628 11047
rect 1618 10961 1628 11017
rect 104 10931 130 10961
rect 1580 10931 1628 10961
rect 1618 10875 1628 10931
rect 104 10845 130 10875
rect 1580 10845 1628 10875
rect 1618 10789 1628 10845
rect 104 10759 130 10789
rect 1580 10759 1628 10789
rect 1618 10703 1628 10759
rect 104 10673 130 10703
rect 1580 10673 1628 10703
rect 1618 10617 1628 10673
rect 104 10587 130 10617
rect 1580 10587 1628 10617
rect 1618 10531 1628 10587
rect 104 10501 130 10531
rect 1580 10501 1628 10531
rect 1618 10445 1628 10501
rect 104 10415 130 10445
rect 1580 10415 1628 10445
rect 1618 10359 1628 10415
rect 104 10329 130 10359
rect 1580 10329 1628 10359
rect 1618 10273 1628 10329
rect 104 10243 130 10273
rect 1580 10243 1628 10273
rect 1618 10187 1628 10243
rect 104 10157 130 10187
rect 1580 10157 1628 10187
rect 1618 10101 1628 10157
rect 104 10071 130 10101
rect 1580 10071 1628 10101
rect 1618 10015 1628 10071
rect 104 9985 130 10015
rect 1580 9985 1628 10015
rect 1618 9929 1628 9985
rect 104 9899 130 9929
rect 1580 9899 1628 9929
rect 1618 9843 1628 9899
rect 104 9813 130 9843
rect 1580 9813 1628 9843
rect 1618 9757 1628 9813
rect 104 9727 130 9757
rect 1580 9727 1628 9757
rect 1618 9671 1628 9727
rect 104 9641 130 9671
rect 1580 9641 1628 9671
rect 1618 9585 1628 9641
rect 104 9555 130 9585
rect 1580 9555 1628 9585
rect 1618 9499 1628 9555
rect 104 9469 130 9499
rect 1580 9469 1628 9499
rect 1618 9413 1628 9469
rect 104 9383 130 9413
rect 1580 9383 1628 9413
rect 1618 9327 1628 9383
rect 104 9297 130 9327
rect 1580 9297 1628 9327
rect 1618 9241 1628 9297
rect 104 9211 130 9241
rect 1580 9211 1628 9241
rect 1618 9155 1628 9211
rect 104 9125 130 9155
rect 1580 9125 1628 9155
rect 1618 9069 1628 9125
rect 104 9039 130 9069
rect 1580 9039 1628 9069
rect 1618 8983 1628 9039
rect 104 8953 130 8983
rect 1580 8953 1628 8983
rect 1618 8897 1628 8953
rect 104 8867 130 8897
rect 1580 8867 1628 8897
rect 1618 8811 1628 8867
rect 104 8781 130 8811
rect 1580 8781 1628 8811
rect 1618 8725 1628 8781
rect 104 8695 130 8725
rect 1580 8695 1628 8725
rect 1618 8639 1628 8695
rect 104 8609 130 8639
rect 1580 8609 1628 8639
rect 1618 8553 1628 8609
rect 104 8523 130 8553
rect 1580 8523 1628 8553
rect 1618 8467 1628 8523
rect 104 8437 130 8467
rect 1580 8437 1628 8467
rect 1618 8381 1628 8437
rect 104 8351 130 8381
rect 1580 8351 1628 8381
rect 1618 8295 1628 8351
rect 104 8265 130 8295
rect 1580 8265 1628 8295
rect 1618 8209 1628 8265
rect 104 8179 130 8209
rect 1580 8179 1628 8209
rect 1618 8123 1628 8179
rect 104 8093 130 8123
rect 1580 8093 1628 8123
rect 1618 8037 1628 8093
rect 104 8007 130 8037
rect 1580 8007 1628 8037
rect 1618 7951 1628 8007
rect 104 7921 130 7951
rect 1580 7921 1628 7951
rect 1618 7865 1628 7921
rect 104 7835 130 7865
rect 1580 7835 1628 7865
rect 1618 7779 1628 7835
rect 104 7749 130 7779
rect 1580 7749 1628 7779
rect 1618 7693 1628 7749
rect 104 7663 130 7693
rect 1580 7663 1628 7693
rect 1618 7607 1628 7663
rect 104 7577 130 7607
rect 1580 7577 1628 7607
rect 1618 7521 1628 7577
rect 104 7491 130 7521
rect 1580 7491 1628 7521
rect 1618 7435 1628 7491
rect 104 7405 130 7435
rect 1580 7405 1628 7435
rect 1618 7349 1628 7405
rect 104 7319 130 7349
rect 1580 7319 1628 7349
rect 1618 7263 1628 7319
rect 104 7233 130 7263
rect 1580 7233 1628 7263
rect 1618 7177 1628 7233
rect 104 7147 130 7177
rect 1580 7147 1628 7177
rect 1618 7091 1628 7147
rect 104 7061 130 7091
rect 1580 7061 1628 7091
rect 1618 7005 1628 7061
rect 104 6975 130 7005
rect 1580 6975 1628 7005
rect 1618 6919 1628 6975
rect 104 6889 130 6919
rect 1580 6889 1628 6919
rect 1618 6833 1628 6889
rect 104 6803 130 6833
rect 1580 6803 1628 6833
rect 1618 6747 1628 6803
rect 104 6717 130 6747
rect 1580 6717 1628 6747
rect 1618 6661 1628 6717
rect 104 6631 130 6661
rect 1580 6631 1628 6661
rect 1618 6575 1628 6631
rect 104 6545 130 6575
rect 1580 6545 1628 6575
rect 1618 6489 1628 6545
rect 104 6459 130 6489
rect 1580 6459 1628 6489
rect 1618 6403 1628 6459
rect 104 6373 130 6403
rect 1580 6373 1628 6403
rect 1618 6317 1628 6373
rect 104 6287 130 6317
rect 1580 6287 1628 6317
rect 1618 6231 1628 6287
rect 104 6201 130 6231
rect 1580 6201 1628 6231
rect 1618 6145 1628 6201
rect 104 6115 130 6145
rect 1580 6115 1628 6145
rect 1618 6059 1628 6115
rect 104 6029 130 6059
rect 1580 6029 1628 6059
rect 1618 5973 1628 6029
rect 104 5943 130 5973
rect 1580 5943 1628 5973
rect 1618 5887 1628 5943
rect 104 5857 130 5887
rect 1580 5857 1628 5887
rect 1618 5801 1628 5857
rect 104 5771 130 5801
rect 1580 5771 1628 5801
rect 1618 5715 1628 5771
rect 104 5685 130 5715
rect 1580 5685 1628 5715
rect 1618 5629 1628 5685
rect 104 5599 130 5629
rect 1580 5599 1628 5629
rect 1618 5543 1628 5599
rect 104 5513 130 5543
rect 1580 5513 1628 5543
rect 1618 5457 1628 5513
rect 104 5427 130 5457
rect 1580 5427 1628 5457
rect 1618 5371 1628 5427
rect 104 5341 130 5371
rect 1580 5341 1628 5371
rect 1618 5285 1628 5341
rect 104 5255 130 5285
rect 1580 5255 1628 5285
rect 1618 5199 1628 5255
rect 104 5169 130 5199
rect 1580 5169 1628 5199
rect 1618 5113 1628 5169
rect 104 5083 130 5113
rect 1580 5083 1628 5113
rect 1618 5027 1628 5083
rect 104 4997 130 5027
rect 1580 4997 1628 5027
rect 1618 4941 1628 4997
rect 104 4911 130 4941
rect 1580 4911 1628 4941
rect 1618 4855 1628 4911
rect 104 4825 130 4855
rect 1580 4825 1628 4855
rect 1618 4769 1628 4825
rect 104 4739 130 4769
rect 1580 4739 1628 4769
rect 1618 4683 1628 4739
rect 104 4653 130 4683
rect 1580 4653 1628 4683
rect 1618 4597 1628 4653
rect 104 4567 130 4597
rect 1580 4567 1628 4597
rect 1618 4511 1628 4567
rect 104 4481 130 4511
rect 1580 4481 1628 4511
rect 1618 4425 1628 4481
rect 104 4395 130 4425
rect 1580 4395 1628 4425
rect 1618 4339 1628 4395
rect 104 4309 130 4339
rect 1580 4309 1628 4339
rect 1618 4253 1628 4309
rect 104 4223 130 4253
rect 1580 4223 1628 4253
rect 1618 4167 1628 4223
rect 104 4137 130 4167
rect 1580 4137 1628 4167
rect 1618 4081 1628 4137
rect 104 4051 130 4081
rect 1580 4051 1628 4081
rect 1618 3995 1628 4051
rect 104 3965 130 3995
rect 1580 3965 1628 3995
rect 1618 3909 1628 3965
rect 104 3879 130 3909
rect 1580 3879 1628 3909
rect 1618 3823 1628 3879
rect 104 3793 130 3823
rect 1580 3793 1628 3823
rect 1618 3737 1628 3793
rect 104 3707 130 3737
rect 1580 3707 1628 3737
rect 1618 3651 1628 3707
rect 104 3621 130 3651
rect 1580 3621 1628 3651
rect 1618 3565 1628 3621
rect 104 3535 130 3565
rect 1580 3535 1628 3565
rect 1618 3479 1628 3535
rect 104 3449 130 3479
rect 1580 3449 1628 3479
rect 1618 3393 1628 3449
rect 104 3363 130 3393
rect 1580 3363 1628 3393
rect 1618 3307 1628 3363
rect 104 3277 130 3307
rect 1580 3277 1628 3307
rect 1618 3221 1628 3277
rect 104 3191 130 3221
rect 1580 3191 1628 3221
rect 1618 3135 1628 3191
rect 104 3105 130 3135
rect 1580 3105 1628 3135
rect 1618 3049 1628 3105
rect 104 3019 130 3049
rect 1580 3019 1628 3049
rect 1618 2963 1628 3019
rect 104 2933 130 2963
rect 1580 2933 1628 2963
rect 1618 2877 1628 2933
rect 104 2847 130 2877
rect 1580 2847 1628 2877
rect 1618 2791 1628 2847
rect 104 2761 130 2791
rect 1580 2761 1628 2791
rect 1618 2705 1628 2761
rect 104 2675 130 2705
rect 1580 2675 1628 2705
rect 1618 2619 1628 2675
rect 104 2589 130 2619
rect 1580 2589 1628 2619
rect 1618 2533 1628 2589
rect 104 2503 130 2533
rect 1580 2503 1628 2533
rect 1618 2447 1628 2503
rect 104 2417 130 2447
rect 1580 2417 1628 2447
rect 1618 2361 1628 2417
rect 104 2331 130 2361
rect 1580 2331 1628 2361
rect 1618 2275 1628 2331
rect 104 2245 130 2275
rect 1580 2245 1628 2275
rect 1618 2189 1628 2245
rect 104 2159 130 2189
rect 1580 2159 1628 2189
rect 1618 2103 1628 2159
rect 104 2073 130 2103
rect 1580 2073 1628 2103
rect 1618 2017 1628 2073
rect 104 1987 130 2017
rect 1580 1987 1628 2017
rect 1618 1931 1628 1987
rect 104 1901 130 1931
rect 1580 1901 1628 1931
rect 1618 1845 1628 1901
rect 104 1815 130 1845
rect 1580 1815 1628 1845
rect 1618 1759 1628 1815
rect 104 1729 130 1759
rect 1580 1729 1628 1759
rect 1618 1673 1628 1729
rect 104 1643 130 1673
rect 1580 1643 1628 1673
rect 1618 1587 1628 1643
rect 104 1557 130 1587
rect 1580 1557 1628 1587
rect 1618 1501 1628 1557
rect 104 1471 130 1501
rect 1580 1471 1628 1501
rect 1618 1415 1628 1471
rect 104 1385 130 1415
rect 1580 1385 1628 1415
rect 1618 1329 1628 1385
rect 104 1299 130 1329
rect 1580 1299 1628 1329
rect 1618 1243 1628 1299
rect 104 1213 130 1243
rect 1580 1213 1628 1243
rect 1618 1157 1628 1213
rect 104 1127 130 1157
rect 1580 1127 1628 1157
rect 1618 1071 1628 1127
rect 104 1041 130 1071
rect 1580 1041 1628 1071
rect 1618 985 1628 1041
rect 104 955 130 985
rect 1580 955 1628 985
rect 1618 899 1628 955
rect 104 869 130 899
rect 1580 869 1628 899
rect 1618 813 1628 869
rect 104 783 130 813
rect 1580 783 1628 813
rect 1618 727 1628 783
rect 104 697 130 727
rect 1580 697 1628 727
rect 1618 641 1628 697
rect 104 611 130 641
rect 1580 611 1628 641
rect 1618 555 1628 611
rect 104 525 130 555
rect 1580 525 1628 555
rect 1618 469 1628 525
rect 104 439 130 469
rect 1580 439 1628 469
rect 1618 383 1628 439
rect 104 353 130 383
rect 1580 353 1628 383
rect 1618 297 1628 353
rect 104 267 130 297
rect 1580 267 1628 297
rect 1618 211 1628 267
rect 104 181 130 211
rect 1580 181 1628 211
rect 1618 179 1628 181
rect 1662 179 1672 43815
rect 1618 163 1672 179
<< polycont >>
rect 1628 179 1662 43815
<< locali >>
rect 36 43924 100 43958
rect 1680 43924 1744 43958
rect 36 43894 70 43924
rect 1710 43894 1744 43924
rect 122 43824 138 43858
rect 1572 43824 1588 43858
rect 1628 43815 1662 43831
rect 122 43738 138 43772
rect 1572 43738 1588 43772
rect 122 43652 138 43686
rect 1572 43652 1588 43686
rect 122 43566 138 43600
rect 1572 43566 1588 43600
rect 122 43480 138 43514
rect 1572 43480 1588 43514
rect 122 43394 138 43428
rect 1572 43394 1588 43428
rect 122 43308 138 43342
rect 1572 43308 1588 43342
rect 122 43222 138 43256
rect 1572 43222 1588 43256
rect 122 43136 138 43170
rect 1572 43136 1588 43170
rect 122 43050 138 43084
rect 1572 43050 1588 43084
rect 122 42964 138 42998
rect 1572 42964 1588 42998
rect 122 42878 138 42912
rect 1572 42878 1588 42912
rect 122 42792 138 42826
rect 1572 42792 1588 42826
rect 122 42706 138 42740
rect 1572 42706 1588 42740
rect 122 42620 138 42654
rect 1572 42620 1588 42654
rect 122 42534 138 42568
rect 1572 42534 1588 42568
rect 122 42448 138 42482
rect 1572 42448 1588 42482
rect 122 42362 138 42396
rect 1572 42362 1588 42396
rect 122 42276 138 42310
rect 1572 42276 1588 42310
rect 122 42190 138 42224
rect 1572 42190 1588 42224
rect 122 42104 138 42138
rect 1572 42104 1588 42138
rect 122 42018 138 42052
rect 1572 42018 1588 42052
rect 122 41932 138 41966
rect 1572 41932 1588 41966
rect 122 41846 138 41880
rect 1572 41846 1588 41880
rect 122 41760 138 41794
rect 1572 41760 1588 41794
rect 122 41674 138 41708
rect 1572 41674 1588 41708
rect 122 41588 138 41622
rect 1572 41588 1588 41622
rect 122 41502 138 41536
rect 1572 41502 1588 41536
rect 122 41416 138 41450
rect 1572 41416 1588 41450
rect 122 41330 138 41364
rect 1572 41330 1588 41364
rect 122 41244 138 41278
rect 1572 41244 1588 41278
rect 122 41158 138 41192
rect 1572 41158 1588 41192
rect 122 41072 138 41106
rect 1572 41072 1588 41106
rect 122 40986 138 41020
rect 1572 40986 1588 41020
rect 122 40900 138 40934
rect 1572 40900 1588 40934
rect 122 40814 138 40848
rect 1572 40814 1588 40848
rect 122 40728 138 40762
rect 1572 40728 1588 40762
rect 122 40642 138 40676
rect 1572 40642 1588 40676
rect 122 40556 138 40590
rect 1572 40556 1588 40590
rect 122 40470 138 40504
rect 1572 40470 1588 40504
rect 122 40384 138 40418
rect 1572 40384 1588 40418
rect 122 40298 138 40332
rect 1572 40298 1588 40332
rect 122 40212 138 40246
rect 1572 40212 1588 40246
rect 122 40126 138 40160
rect 1572 40126 1588 40160
rect 122 40040 138 40074
rect 1572 40040 1588 40074
rect 122 39954 138 39988
rect 1572 39954 1588 39988
rect 122 39868 138 39902
rect 1572 39868 1588 39902
rect 122 39782 138 39816
rect 1572 39782 1588 39816
rect 122 39696 138 39730
rect 1572 39696 1588 39730
rect 122 39610 138 39644
rect 1572 39610 1588 39644
rect 122 39524 138 39558
rect 1572 39524 1588 39558
rect 122 39438 138 39472
rect 1572 39438 1588 39472
rect 122 39352 138 39386
rect 1572 39352 1588 39386
rect 122 39266 138 39300
rect 1572 39266 1588 39300
rect 122 39180 138 39214
rect 1572 39180 1588 39214
rect 122 39094 138 39128
rect 1572 39094 1588 39128
rect 122 39008 138 39042
rect 1572 39008 1588 39042
rect 122 38922 138 38956
rect 1572 38922 1588 38956
rect 122 38836 138 38870
rect 1572 38836 1588 38870
rect 122 38750 138 38784
rect 1572 38750 1588 38784
rect 122 38664 138 38698
rect 1572 38664 1588 38698
rect 122 38578 138 38612
rect 1572 38578 1588 38612
rect 122 38492 138 38526
rect 1572 38492 1588 38526
rect 122 38406 138 38440
rect 1572 38406 1588 38440
rect 122 38320 138 38354
rect 1572 38320 1588 38354
rect 122 38234 138 38268
rect 1572 38234 1588 38268
rect 122 38148 138 38182
rect 1572 38148 1588 38182
rect 122 38062 138 38096
rect 1572 38062 1588 38096
rect 122 37976 138 38010
rect 1572 37976 1588 38010
rect 122 37890 138 37924
rect 1572 37890 1588 37924
rect 122 37804 138 37838
rect 1572 37804 1588 37838
rect 122 37718 138 37752
rect 1572 37718 1588 37752
rect 122 37632 138 37666
rect 1572 37632 1588 37666
rect 122 37546 138 37580
rect 1572 37546 1588 37580
rect 122 37460 138 37494
rect 1572 37460 1588 37494
rect 122 37374 138 37408
rect 1572 37374 1588 37408
rect 122 37288 138 37322
rect 1572 37288 1588 37322
rect 122 37202 138 37236
rect 1572 37202 1588 37236
rect 122 37116 138 37150
rect 1572 37116 1588 37150
rect 122 37030 138 37064
rect 1572 37030 1588 37064
rect 122 36944 138 36978
rect 1572 36944 1588 36978
rect 122 36858 138 36892
rect 1572 36858 1588 36892
rect 122 36772 138 36806
rect 1572 36772 1588 36806
rect 122 36686 138 36720
rect 1572 36686 1588 36720
rect 122 36600 138 36634
rect 1572 36600 1588 36634
rect 122 36514 138 36548
rect 1572 36514 1588 36548
rect 122 36428 138 36462
rect 1572 36428 1588 36462
rect 122 36342 138 36376
rect 1572 36342 1588 36376
rect 122 36256 138 36290
rect 1572 36256 1588 36290
rect 122 36170 138 36204
rect 1572 36170 1588 36204
rect 122 36084 138 36118
rect 1572 36084 1588 36118
rect 122 35998 138 36032
rect 1572 35998 1588 36032
rect 122 35912 138 35946
rect 1572 35912 1588 35946
rect 122 35826 138 35860
rect 1572 35826 1588 35860
rect 122 35740 138 35774
rect 1572 35740 1588 35774
rect 122 35654 138 35688
rect 1572 35654 1588 35688
rect 122 35568 138 35602
rect 1572 35568 1588 35602
rect 122 35482 138 35516
rect 1572 35482 1588 35516
rect 122 35396 138 35430
rect 1572 35396 1588 35430
rect 122 35310 138 35344
rect 1572 35310 1588 35344
rect 122 35224 138 35258
rect 1572 35224 1588 35258
rect 122 35138 138 35172
rect 1572 35138 1588 35172
rect 122 35052 138 35086
rect 1572 35052 1588 35086
rect 122 34966 138 35000
rect 1572 34966 1588 35000
rect 122 34880 138 34914
rect 1572 34880 1588 34914
rect 122 34794 138 34828
rect 1572 34794 1588 34828
rect 122 34708 138 34742
rect 1572 34708 1588 34742
rect 122 34622 138 34656
rect 1572 34622 1588 34656
rect 122 34536 138 34570
rect 1572 34536 1588 34570
rect 122 34450 138 34484
rect 1572 34450 1588 34484
rect 122 34364 138 34398
rect 1572 34364 1588 34398
rect 122 34278 138 34312
rect 1572 34278 1588 34312
rect 122 34192 138 34226
rect 1572 34192 1588 34226
rect 122 34106 138 34140
rect 1572 34106 1588 34140
rect 122 34020 138 34054
rect 1572 34020 1588 34054
rect 122 33934 138 33968
rect 1572 33934 1588 33968
rect 122 33848 138 33882
rect 1572 33848 1588 33882
rect 122 33762 138 33796
rect 1572 33762 1588 33796
rect 122 33676 138 33710
rect 1572 33676 1588 33710
rect 122 33590 138 33624
rect 1572 33590 1588 33624
rect 122 33504 138 33538
rect 1572 33504 1588 33538
rect 122 33418 138 33452
rect 1572 33418 1588 33452
rect 122 33332 138 33366
rect 1572 33332 1588 33366
rect 122 33246 138 33280
rect 1572 33246 1588 33280
rect 122 33160 138 33194
rect 1572 33160 1588 33194
rect 122 33074 138 33108
rect 1572 33074 1588 33108
rect 122 32988 138 33022
rect 1572 32988 1588 33022
rect 122 32902 138 32936
rect 1572 32902 1588 32936
rect 122 32816 138 32850
rect 1572 32816 1588 32850
rect 122 32730 138 32764
rect 1572 32730 1588 32764
rect 122 32644 138 32678
rect 1572 32644 1588 32678
rect 122 32558 138 32592
rect 1572 32558 1588 32592
rect 122 32472 138 32506
rect 1572 32472 1588 32506
rect 122 32386 138 32420
rect 1572 32386 1588 32420
rect 122 32300 138 32334
rect 1572 32300 1588 32334
rect 122 32214 138 32248
rect 1572 32214 1588 32248
rect 122 32128 138 32162
rect 1572 32128 1588 32162
rect 122 32042 138 32076
rect 1572 32042 1588 32076
rect 122 31956 138 31990
rect 1572 31956 1588 31990
rect 122 31870 138 31904
rect 1572 31870 1588 31904
rect 122 31784 138 31818
rect 1572 31784 1588 31818
rect 122 31698 138 31732
rect 1572 31698 1588 31732
rect 122 31612 138 31646
rect 1572 31612 1588 31646
rect 122 31526 138 31560
rect 1572 31526 1588 31560
rect 122 31440 138 31474
rect 1572 31440 1588 31474
rect 122 31354 138 31388
rect 1572 31354 1588 31388
rect 122 31268 138 31302
rect 1572 31268 1588 31302
rect 122 31182 138 31216
rect 1572 31182 1588 31216
rect 122 31096 138 31130
rect 1572 31096 1588 31130
rect 122 31010 138 31044
rect 1572 31010 1588 31044
rect 122 30924 138 30958
rect 1572 30924 1588 30958
rect 122 30838 138 30872
rect 1572 30838 1588 30872
rect 122 30752 138 30786
rect 1572 30752 1588 30786
rect 122 30666 138 30700
rect 1572 30666 1588 30700
rect 122 30580 138 30614
rect 1572 30580 1588 30614
rect 122 30494 138 30528
rect 1572 30494 1588 30528
rect 122 30408 138 30442
rect 1572 30408 1588 30442
rect 122 30322 138 30356
rect 1572 30322 1588 30356
rect 122 30236 138 30270
rect 1572 30236 1588 30270
rect 122 30150 138 30184
rect 1572 30150 1588 30184
rect 122 30064 138 30098
rect 1572 30064 1588 30098
rect 122 29978 138 30012
rect 1572 29978 1588 30012
rect 122 29892 138 29926
rect 1572 29892 1588 29926
rect 122 29806 138 29840
rect 1572 29806 1588 29840
rect 122 29720 138 29754
rect 1572 29720 1588 29754
rect 122 29634 138 29668
rect 1572 29634 1588 29668
rect 122 29548 138 29582
rect 1572 29548 1588 29582
rect 122 29462 138 29496
rect 1572 29462 1588 29496
rect 122 29376 138 29410
rect 1572 29376 1588 29410
rect 122 29290 138 29324
rect 1572 29290 1588 29324
rect 122 29204 138 29238
rect 1572 29204 1588 29238
rect 122 29118 138 29152
rect 1572 29118 1588 29152
rect 122 29032 138 29066
rect 1572 29032 1588 29066
rect 122 28946 138 28980
rect 1572 28946 1588 28980
rect 122 28860 138 28894
rect 1572 28860 1588 28894
rect 122 28774 138 28808
rect 1572 28774 1588 28808
rect 122 28688 138 28722
rect 1572 28688 1588 28722
rect 122 28602 138 28636
rect 1572 28602 1588 28636
rect 122 28516 138 28550
rect 1572 28516 1588 28550
rect 122 28430 138 28464
rect 1572 28430 1588 28464
rect 122 28344 138 28378
rect 1572 28344 1588 28378
rect 122 28258 138 28292
rect 1572 28258 1588 28292
rect 122 28172 138 28206
rect 1572 28172 1588 28206
rect 122 28086 138 28120
rect 1572 28086 1588 28120
rect 122 28000 138 28034
rect 1572 28000 1588 28034
rect 122 27914 138 27948
rect 1572 27914 1588 27948
rect 122 27828 138 27862
rect 1572 27828 1588 27862
rect 122 27742 138 27776
rect 1572 27742 1588 27776
rect 122 27656 138 27690
rect 1572 27656 1588 27690
rect 122 27570 138 27604
rect 1572 27570 1588 27604
rect 122 27484 138 27518
rect 1572 27484 1588 27518
rect 122 27398 138 27432
rect 1572 27398 1588 27432
rect 122 27312 138 27346
rect 1572 27312 1588 27346
rect 122 27226 138 27260
rect 1572 27226 1588 27260
rect 122 27140 138 27174
rect 1572 27140 1588 27174
rect 122 27054 138 27088
rect 1572 27054 1588 27088
rect 122 26968 138 27002
rect 1572 26968 1588 27002
rect 122 26882 138 26916
rect 1572 26882 1588 26916
rect 122 26796 138 26830
rect 1572 26796 1588 26830
rect 122 26710 138 26744
rect 1572 26710 1588 26744
rect 122 26624 138 26658
rect 1572 26624 1588 26658
rect 122 26538 138 26572
rect 1572 26538 1588 26572
rect 122 26452 138 26486
rect 1572 26452 1588 26486
rect 122 26366 138 26400
rect 1572 26366 1588 26400
rect 122 26280 138 26314
rect 1572 26280 1588 26314
rect 122 26194 138 26228
rect 1572 26194 1588 26228
rect 122 26108 138 26142
rect 1572 26108 1588 26142
rect 122 26022 138 26056
rect 1572 26022 1588 26056
rect 122 25936 138 25970
rect 1572 25936 1588 25970
rect 122 25850 138 25884
rect 1572 25850 1588 25884
rect 122 25764 138 25798
rect 1572 25764 1588 25798
rect 122 25678 138 25712
rect 1572 25678 1588 25712
rect 122 25592 138 25626
rect 1572 25592 1588 25626
rect 122 25506 138 25540
rect 1572 25506 1588 25540
rect 122 25420 138 25454
rect 1572 25420 1588 25454
rect 122 25334 138 25368
rect 1572 25334 1588 25368
rect 122 25248 138 25282
rect 1572 25248 1588 25282
rect 122 25162 138 25196
rect 1572 25162 1588 25196
rect 122 25076 138 25110
rect 1572 25076 1588 25110
rect 122 24990 138 25024
rect 1572 24990 1588 25024
rect 122 24904 138 24938
rect 1572 24904 1588 24938
rect 122 24818 138 24852
rect 1572 24818 1588 24852
rect 122 24732 138 24766
rect 1572 24732 1588 24766
rect 122 24646 138 24680
rect 1572 24646 1588 24680
rect 122 24560 138 24594
rect 1572 24560 1588 24594
rect 122 24474 138 24508
rect 1572 24474 1588 24508
rect 122 24388 138 24422
rect 1572 24388 1588 24422
rect 122 24302 138 24336
rect 1572 24302 1588 24336
rect 122 24216 138 24250
rect 1572 24216 1588 24250
rect 122 24130 138 24164
rect 1572 24130 1588 24164
rect 122 24044 138 24078
rect 1572 24044 1588 24078
rect 122 23958 138 23992
rect 1572 23958 1588 23992
rect 122 23872 138 23906
rect 1572 23872 1588 23906
rect 122 23786 138 23820
rect 1572 23786 1588 23820
rect 122 23700 138 23734
rect 1572 23700 1588 23734
rect 122 23614 138 23648
rect 1572 23614 1588 23648
rect 122 23528 138 23562
rect 1572 23528 1588 23562
rect 122 23442 138 23476
rect 1572 23442 1588 23476
rect 122 23356 138 23390
rect 1572 23356 1588 23390
rect 122 23270 138 23304
rect 1572 23270 1588 23304
rect 122 23184 138 23218
rect 1572 23184 1588 23218
rect 122 23098 138 23132
rect 1572 23098 1588 23132
rect 122 23012 138 23046
rect 1572 23012 1588 23046
rect 122 22926 138 22960
rect 1572 22926 1588 22960
rect 122 22840 138 22874
rect 1572 22840 1588 22874
rect 122 22754 138 22788
rect 1572 22754 1588 22788
rect 122 22668 138 22702
rect 1572 22668 1588 22702
rect 122 22582 138 22616
rect 1572 22582 1588 22616
rect 122 22496 138 22530
rect 1572 22496 1588 22530
rect 122 22410 138 22444
rect 1572 22410 1588 22444
rect 122 22324 138 22358
rect 1572 22324 1588 22358
rect 122 22238 138 22272
rect 1572 22238 1588 22272
rect 122 22152 138 22186
rect 1572 22152 1588 22186
rect 122 22066 138 22100
rect 1572 22066 1588 22100
rect 122 21980 138 22014
rect 1572 21980 1588 22014
rect 122 21894 138 21928
rect 1572 21894 1588 21928
rect 122 21808 138 21842
rect 1572 21808 1588 21842
rect 122 21722 138 21756
rect 1572 21722 1588 21756
rect 122 21636 138 21670
rect 1572 21636 1588 21670
rect 122 21550 138 21584
rect 1572 21550 1588 21584
rect 122 21464 138 21498
rect 1572 21464 1588 21498
rect 122 21378 138 21412
rect 1572 21378 1588 21412
rect 122 21292 138 21326
rect 1572 21292 1588 21326
rect 122 21206 138 21240
rect 1572 21206 1588 21240
rect 122 21120 138 21154
rect 1572 21120 1588 21154
rect 122 21034 138 21068
rect 1572 21034 1588 21068
rect 122 20948 138 20982
rect 1572 20948 1588 20982
rect 122 20862 138 20896
rect 1572 20862 1588 20896
rect 122 20776 138 20810
rect 1572 20776 1588 20810
rect 122 20690 138 20724
rect 1572 20690 1588 20724
rect 122 20604 138 20638
rect 1572 20604 1588 20638
rect 122 20518 138 20552
rect 1572 20518 1588 20552
rect 122 20432 138 20466
rect 1572 20432 1588 20466
rect 122 20346 138 20380
rect 1572 20346 1588 20380
rect 122 20260 138 20294
rect 1572 20260 1588 20294
rect 122 20174 138 20208
rect 1572 20174 1588 20208
rect 122 20088 138 20122
rect 1572 20088 1588 20122
rect 122 20002 138 20036
rect 1572 20002 1588 20036
rect 122 19916 138 19950
rect 1572 19916 1588 19950
rect 122 19830 138 19864
rect 1572 19830 1588 19864
rect 122 19744 138 19778
rect 1572 19744 1588 19778
rect 122 19658 138 19692
rect 1572 19658 1588 19692
rect 122 19572 138 19606
rect 1572 19572 1588 19606
rect 122 19486 138 19520
rect 1572 19486 1588 19520
rect 122 19400 138 19434
rect 1572 19400 1588 19434
rect 122 19314 138 19348
rect 1572 19314 1588 19348
rect 122 19228 138 19262
rect 1572 19228 1588 19262
rect 122 19142 138 19176
rect 1572 19142 1588 19176
rect 122 19056 138 19090
rect 1572 19056 1588 19090
rect 122 18970 138 19004
rect 1572 18970 1588 19004
rect 122 18884 138 18918
rect 1572 18884 1588 18918
rect 122 18798 138 18832
rect 1572 18798 1588 18832
rect 122 18712 138 18746
rect 1572 18712 1588 18746
rect 122 18626 138 18660
rect 1572 18626 1588 18660
rect 122 18540 138 18574
rect 1572 18540 1588 18574
rect 122 18454 138 18488
rect 1572 18454 1588 18488
rect 122 18368 138 18402
rect 1572 18368 1588 18402
rect 122 18282 138 18316
rect 1572 18282 1588 18316
rect 122 18196 138 18230
rect 1572 18196 1588 18230
rect 122 18110 138 18144
rect 1572 18110 1588 18144
rect 122 18024 138 18058
rect 1572 18024 1588 18058
rect 122 17938 138 17972
rect 1572 17938 1588 17972
rect 122 17852 138 17886
rect 1572 17852 1588 17886
rect 122 17766 138 17800
rect 1572 17766 1588 17800
rect 122 17680 138 17714
rect 1572 17680 1588 17714
rect 122 17594 138 17628
rect 1572 17594 1588 17628
rect 122 17508 138 17542
rect 1572 17508 1588 17542
rect 122 17422 138 17456
rect 1572 17422 1588 17456
rect 122 17336 138 17370
rect 1572 17336 1588 17370
rect 122 17250 138 17284
rect 1572 17250 1588 17284
rect 122 17164 138 17198
rect 1572 17164 1588 17198
rect 122 17078 138 17112
rect 1572 17078 1588 17112
rect 122 16992 138 17026
rect 1572 16992 1588 17026
rect 122 16906 138 16940
rect 1572 16906 1588 16940
rect 122 16820 138 16854
rect 1572 16820 1588 16854
rect 122 16734 138 16768
rect 1572 16734 1588 16768
rect 122 16648 138 16682
rect 1572 16648 1588 16682
rect 122 16562 138 16596
rect 1572 16562 1588 16596
rect 122 16476 138 16510
rect 1572 16476 1588 16510
rect 122 16390 138 16424
rect 1572 16390 1588 16424
rect 122 16304 138 16338
rect 1572 16304 1588 16338
rect 122 16218 138 16252
rect 1572 16218 1588 16252
rect 122 16132 138 16166
rect 1572 16132 1588 16166
rect 122 16046 138 16080
rect 1572 16046 1588 16080
rect 122 15960 138 15994
rect 1572 15960 1588 15994
rect 122 15874 138 15908
rect 1572 15874 1588 15908
rect 122 15788 138 15822
rect 1572 15788 1588 15822
rect 122 15702 138 15736
rect 1572 15702 1588 15736
rect 122 15616 138 15650
rect 1572 15616 1588 15650
rect 122 15530 138 15564
rect 1572 15530 1588 15564
rect 122 15444 138 15478
rect 1572 15444 1588 15478
rect 122 15358 138 15392
rect 1572 15358 1588 15392
rect 122 15272 138 15306
rect 1572 15272 1588 15306
rect 122 15186 138 15220
rect 1572 15186 1588 15220
rect 122 15100 138 15134
rect 1572 15100 1588 15134
rect 122 15014 138 15048
rect 1572 15014 1588 15048
rect 122 14928 138 14962
rect 1572 14928 1588 14962
rect 122 14842 138 14876
rect 1572 14842 1588 14876
rect 122 14756 138 14790
rect 1572 14756 1588 14790
rect 122 14670 138 14704
rect 1572 14670 1588 14704
rect 122 14584 138 14618
rect 1572 14584 1588 14618
rect 122 14498 138 14532
rect 1572 14498 1588 14532
rect 122 14412 138 14446
rect 1572 14412 1588 14446
rect 122 14326 138 14360
rect 1572 14326 1588 14360
rect 122 14240 138 14274
rect 1572 14240 1588 14274
rect 122 14154 138 14188
rect 1572 14154 1588 14188
rect 122 14068 138 14102
rect 1572 14068 1588 14102
rect 122 13982 138 14016
rect 1572 13982 1588 14016
rect 122 13896 138 13930
rect 1572 13896 1588 13930
rect 122 13810 138 13844
rect 1572 13810 1588 13844
rect 122 13724 138 13758
rect 1572 13724 1588 13758
rect 122 13638 138 13672
rect 1572 13638 1588 13672
rect 122 13552 138 13586
rect 1572 13552 1588 13586
rect 122 13466 138 13500
rect 1572 13466 1588 13500
rect 122 13380 138 13414
rect 1572 13380 1588 13414
rect 122 13294 138 13328
rect 1572 13294 1588 13328
rect 122 13208 138 13242
rect 1572 13208 1588 13242
rect 122 13122 138 13156
rect 1572 13122 1588 13156
rect 122 13036 138 13070
rect 1572 13036 1588 13070
rect 122 12950 138 12984
rect 1572 12950 1588 12984
rect 122 12864 138 12898
rect 1572 12864 1588 12898
rect 122 12778 138 12812
rect 1572 12778 1588 12812
rect 122 12692 138 12726
rect 1572 12692 1588 12726
rect 122 12606 138 12640
rect 1572 12606 1588 12640
rect 122 12520 138 12554
rect 1572 12520 1588 12554
rect 122 12434 138 12468
rect 1572 12434 1588 12468
rect 122 12348 138 12382
rect 1572 12348 1588 12382
rect 122 12262 138 12296
rect 1572 12262 1588 12296
rect 122 12176 138 12210
rect 1572 12176 1588 12210
rect 122 12090 138 12124
rect 1572 12090 1588 12124
rect 122 12004 138 12038
rect 1572 12004 1588 12038
rect 122 11918 138 11952
rect 1572 11918 1588 11952
rect 122 11832 138 11866
rect 1572 11832 1588 11866
rect 122 11746 138 11780
rect 1572 11746 1588 11780
rect 122 11660 138 11694
rect 1572 11660 1588 11694
rect 122 11574 138 11608
rect 1572 11574 1588 11608
rect 122 11488 138 11522
rect 1572 11488 1588 11522
rect 122 11402 138 11436
rect 1572 11402 1588 11436
rect 122 11316 138 11350
rect 1572 11316 1588 11350
rect 122 11230 138 11264
rect 1572 11230 1588 11264
rect 122 11144 138 11178
rect 1572 11144 1588 11178
rect 122 11058 138 11092
rect 1572 11058 1588 11092
rect 122 10972 138 11006
rect 1572 10972 1588 11006
rect 122 10886 138 10920
rect 1572 10886 1588 10920
rect 122 10800 138 10834
rect 1572 10800 1588 10834
rect 122 10714 138 10748
rect 1572 10714 1588 10748
rect 122 10628 138 10662
rect 1572 10628 1588 10662
rect 122 10542 138 10576
rect 1572 10542 1588 10576
rect 122 10456 138 10490
rect 1572 10456 1588 10490
rect 122 10370 138 10404
rect 1572 10370 1588 10404
rect 122 10284 138 10318
rect 1572 10284 1588 10318
rect 122 10198 138 10232
rect 1572 10198 1588 10232
rect 122 10112 138 10146
rect 1572 10112 1588 10146
rect 122 10026 138 10060
rect 1572 10026 1588 10060
rect 122 9940 138 9974
rect 1572 9940 1588 9974
rect 122 9854 138 9888
rect 1572 9854 1588 9888
rect 122 9768 138 9802
rect 1572 9768 1588 9802
rect 122 9682 138 9716
rect 1572 9682 1588 9716
rect 122 9596 138 9630
rect 1572 9596 1588 9630
rect 122 9510 138 9544
rect 1572 9510 1588 9544
rect 122 9424 138 9458
rect 1572 9424 1588 9458
rect 122 9338 138 9372
rect 1572 9338 1588 9372
rect 122 9252 138 9286
rect 1572 9252 1588 9286
rect 122 9166 138 9200
rect 1572 9166 1588 9200
rect 122 9080 138 9114
rect 1572 9080 1588 9114
rect 122 8994 138 9028
rect 1572 8994 1588 9028
rect 122 8908 138 8942
rect 1572 8908 1588 8942
rect 122 8822 138 8856
rect 1572 8822 1588 8856
rect 122 8736 138 8770
rect 1572 8736 1588 8770
rect 122 8650 138 8684
rect 1572 8650 1588 8684
rect 122 8564 138 8598
rect 1572 8564 1588 8598
rect 122 8478 138 8512
rect 1572 8478 1588 8512
rect 122 8392 138 8426
rect 1572 8392 1588 8426
rect 122 8306 138 8340
rect 1572 8306 1588 8340
rect 122 8220 138 8254
rect 1572 8220 1588 8254
rect 122 8134 138 8168
rect 1572 8134 1588 8168
rect 122 8048 138 8082
rect 1572 8048 1588 8082
rect 122 7962 138 7996
rect 1572 7962 1588 7996
rect 122 7876 138 7910
rect 1572 7876 1588 7910
rect 122 7790 138 7824
rect 1572 7790 1588 7824
rect 122 7704 138 7738
rect 1572 7704 1588 7738
rect 122 7618 138 7652
rect 1572 7618 1588 7652
rect 122 7532 138 7566
rect 1572 7532 1588 7566
rect 122 7446 138 7480
rect 1572 7446 1588 7480
rect 122 7360 138 7394
rect 1572 7360 1588 7394
rect 122 7274 138 7308
rect 1572 7274 1588 7308
rect 122 7188 138 7222
rect 1572 7188 1588 7222
rect 122 7102 138 7136
rect 1572 7102 1588 7136
rect 122 7016 138 7050
rect 1572 7016 1588 7050
rect 122 6930 138 6964
rect 1572 6930 1588 6964
rect 122 6844 138 6878
rect 1572 6844 1588 6878
rect 122 6758 138 6792
rect 1572 6758 1588 6792
rect 122 6672 138 6706
rect 1572 6672 1588 6706
rect 122 6586 138 6620
rect 1572 6586 1588 6620
rect 122 6500 138 6534
rect 1572 6500 1588 6534
rect 122 6414 138 6448
rect 1572 6414 1588 6448
rect 122 6328 138 6362
rect 1572 6328 1588 6362
rect 122 6242 138 6276
rect 1572 6242 1588 6276
rect 122 6156 138 6190
rect 1572 6156 1588 6190
rect 122 6070 138 6104
rect 1572 6070 1588 6104
rect 122 5984 138 6018
rect 1572 5984 1588 6018
rect 122 5898 138 5932
rect 1572 5898 1588 5932
rect 122 5812 138 5846
rect 1572 5812 1588 5846
rect 122 5726 138 5760
rect 1572 5726 1588 5760
rect 122 5640 138 5674
rect 1572 5640 1588 5674
rect 122 5554 138 5588
rect 1572 5554 1588 5588
rect 122 5468 138 5502
rect 1572 5468 1588 5502
rect 122 5382 138 5416
rect 1572 5382 1588 5416
rect 122 5296 138 5330
rect 1572 5296 1588 5330
rect 122 5210 138 5244
rect 1572 5210 1588 5244
rect 122 5124 138 5158
rect 1572 5124 1588 5158
rect 122 5038 138 5072
rect 1572 5038 1588 5072
rect 122 4952 138 4986
rect 1572 4952 1588 4986
rect 122 4866 138 4900
rect 1572 4866 1588 4900
rect 122 4780 138 4814
rect 1572 4780 1588 4814
rect 122 4694 138 4728
rect 1572 4694 1588 4728
rect 122 4608 138 4642
rect 1572 4608 1588 4642
rect 122 4522 138 4556
rect 1572 4522 1588 4556
rect 122 4436 138 4470
rect 1572 4436 1588 4470
rect 122 4350 138 4384
rect 1572 4350 1588 4384
rect 122 4264 138 4298
rect 1572 4264 1588 4298
rect 122 4178 138 4212
rect 1572 4178 1588 4212
rect 122 4092 138 4126
rect 1572 4092 1588 4126
rect 122 4006 138 4040
rect 1572 4006 1588 4040
rect 122 3920 138 3954
rect 1572 3920 1588 3954
rect 122 3834 138 3868
rect 1572 3834 1588 3868
rect 122 3748 138 3782
rect 1572 3748 1588 3782
rect 122 3662 138 3696
rect 1572 3662 1588 3696
rect 122 3576 138 3610
rect 1572 3576 1588 3610
rect 122 3490 138 3524
rect 1572 3490 1588 3524
rect 122 3404 138 3438
rect 1572 3404 1588 3438
rect 122 3318 138 3352
rect 1572 3318 1588 3352
rect 122 3232 138 3266
rect 1572 3232 1588 3266
rect 122 3146 138 3180
rect 1572 3146 1588 3180
rect 122 3060 138 3094
rect 1572 3060 1588 3094
rect 122 2974 138 3008
rect 1572 2974 1588 3008
rect 122 2888 138 2922
rect 1572 2888 1588 2922
rect 122 2802 138 2836
rect 1572 2802 1588 2836
rect 122 2716 138 2750
rect 1572 2716 1588 2750
rect 122 2630 138 2664
rect 1572 2630 1588 2664
rect 122 2544 138 2578
rect 1572 2544 1588 2578
rect 122 2458 138 2492
rect 1572 2458 1588 2492
rect 122 2372 138 2406
rect 1572 2372 1588 2406
rect 122 2286 138 2320
rect 1572 2286 1588 2320
rect 122 2200 138 2234
rect 1572 2200 1588 2234
rect 122 2114 138 2148
rect 1572 2114 1588 2148
rect 122 2028 138 2062
rect 1572 2028 1588 2062
rect 122 1942 138 1976
rect 1572 1942 1588 1976
rect 122 1856 138 1890
rect 1572 1856 1588 1890
rect 122 1770 138 1804
rect 1572 1770 1588 1804
rect 122 1684 138 1718
rect 1572 1684 1588 1718
rect 122 1598 138 1632
rect 1572 1598 1588 1632
rect 122 1512 138 1546
rect 1572 1512 1588 1546
rect 122 1426 138 1460
rect 1572 1426 1588 1460
rect 122 1340 138 1374
rect 1572 1340 1588 1374
rect 122 1254 138 1288
rect 1572 1254 1588 1288
rect 122 1168 138 1202
rect 1572 1168 1588 1202
rect 122 1082 138 1116
rect 1572 1082 1588 1116
rect 122 996 138 1030
rect 1572 996 1588 1030
rect 122 910 138 944
rect 1572 910 1588 944
rect 122 824 138 858
rect 1572 824 1588 858
rect 122 738 138 772
rect 1572 738 1588 772
rect 122 652 138 686
rect 1572 652 1588 686
rect 122 566 138 600
rect 1572 566 1588 600
rect 122 480 138 514
rect 1572 480 1588 514
rect 122 394 138 428
rect 1572 394 1588 428
rect 122 308 138 342
rect 1572 308 1588 342
rect 122 222 138 256
rect 1572 222 1588 256
rect 122 136 138 170
rect 1572 136 1588 170
rect 1628 163 1662 179
rect 36 70 70 100
rect 1710 70 1744 100
rect 36 36 100 70
rect 1680 36 1744 70
<< viali >>
rect 100 43924 1680 43958
rect 36 100 70 43894
rect 138 43824 1572 43858
rect 138 43738 1572 43772
rect 138 43652 1572 43686
rect 138 43566 1572 43600
rect 138 43480 1572 43514
rect 138 43394 1572 43428
rect 138 43308 1572 43342
rect 138 43222 1572 43256
rect 138 43136 1572 43170
rect 138 43050 1572 43084
rect 138 42964 1572 42998
rect 138 42878 1572 42912
rect 138 42792 1572 42826
rect 138 42706 1572 42740
rect 138 42620 1572 42654
rect 138 42534 1572 42568
rect 138 42448 1572 42482
rect 138 42362 1572 42396
rect 138 42276 1572 42310
rect 138 42190 1572 42224
rect 138 42104 1572 42138
rect 138 42018 1572 42052
rect 138 41932 1572 41966
rect 138 41846 1572 41880
rect 138 41760 1572 41794
rect 138 41674 1572 41708
rect 138 41588 1572 41622
rect 138 41502 1572 41536
rect 138 41416 1572 41450
rect 138 41330 1572 41364
rect 138 41244 1572 41278
rect 138 41158 1572 41192
rect 138 41072 1572 41106
rect 138 40986 1572 41020
rect 138 40900 1572 40934
rect 138 40814 1572 40848
rect 138 40728 1572 40762
rect 138 40642 1572 40676
rect 138 40556 1572 40590
rect 138 40470 1572 40504
rect 138 40384 1572 40418
rect 138 40298 1572 40332
rect 138 40212 1572 40246
rect 138 40126 1572 40160
rect 138 40040 1572 40074
rect 138 39954 1572 39988
rect 138 39868 1572 39902
rect 138 39782 1572 39816
rect 138 39696 1572 39730
rect 138 39610 1572 39644
rect 138 39524 1572 39558
rect 138 39438 1572 39472
rect 138 39352 1572 39386
rect 138 39266 1572 39300
rect 138 39180 1572 39214
rect 138 39094 1572 39128
rect 138 39008 1572 39042
rect 138 38922 1572 38956
rect 138 38836 1572 38870
rect 138 38750 1572 38784
rect 138 38664 1572 38698
rect 138 38578 1572 38612
rect 138 38492 1572 38526
rect 138 38406 1572 38440
rect 138 38320 1572 38354
rect 138 38234 1572 38268
rect 138 38148 1572 38182
rect 138 38062 1572 38096
rect 138 37976 1572 38010
rect 138 37890 1572 37924
rect 138 37804 1572 37838
rect 138 37718 1572 37752
rect 138 37632 1572 37666
rect 138 37546 1572 37580
rect 138 37460 1572 37494
rect 138 37374 1572 37408
rect 138 37288 1572 37322
rect 138 37202 1572 37236
rect 138 37116 1572 37150
rect 138 37030 1572 37064
rect 138 36944 1572 36978
rect 138 36858 1572 36892
rect 138 36772 1572 36806
rect 138 36686 1572 36720
rect 138 36600 1572 36634
rect 138 36514 1572 36548
rect 138 36428 1572 36462
rect 138 36342 1572 36376
rect 138 36256 1572 36290
rect 138 36170 1572 36204
rect 138 36084 1572 36118
rect 138 35998 1572 36032
rect 138 35912 1572 35946
rect 138 35826 1572 35860
rect 138 35740 1572 35774
rect 138 35654 1572 35688
rect 138 35568 1572 35602
rect 138 35482 1572 35516
rect 138 35396 1572 35430
rect 138 35310 1572 35344
rect 138 35224 1572 35258
rect 138 35138 1572 35172
rect 138 35052 1572 35086
rect 138 34966 1572 35000
rect 138 34880 1572 34914
rect 138 34794 1572 34828
rect 138 34708 1572 34742
rect 138 34622 1572 34656
rect 138 34536 1572 34570
rect 138 34450 1572 34484
rect 138 34364 1572 34398
rect 138 34278 1572 34312
rect 138 34192 1572 34226
rect 138 34106 1572 34140
rect 138 34020 1572 34054
rect 138 33934 1572 33968
rect 138 33848 1572 33882
rect 138 33762 1572 33796
rect 138 33676 1572 33710
rect 138 33590 1572 33624
rect 138 33504 1572 33538
rect 138 33418 1572 33452
rect 138 33332 1572 33366
rect 138 33246 1572 33280
rect 138 33160 1572 33194
rect 138 33074 1572 33108
rect 138 32988 1572 33022
rect 138 32902 1572 32936
rect 138 32816 1572 32850
rect 138 32730 1572 32764
rect 138 32644 1572 32678
rect 138 32558 1572 32592
rect 138 32472 1572 32506
rect 138 32386 1572 32420
rect 138 32300 1572 32334
rect 138 32214 1572 32248
rect 138 32128 1572 32162
rect 138 32042 1572 32076
rect 138 31956 1572 31990
rect 138 31870 1572 31904
rect 138 31784 1572 31818
rect 138 31698 1572 31732
rect 138 31612 1572 31646
rect 138 31526 1572 31560
rect 138 31440 1572 31474
rect 138 31354 1572 31388
rect 138 31268 1572 31302
rect 138 31182 1572 31216
rect 138 31096 1572 31130
rect 138 31010 1572 31044
rect 138 30924 1572 30958
rect 138 30838 1572 30872
rect 138 30752 1572 30786
rect 138 30666 1572 30700
rect 138 30580 1572 30614
rect 138 30494 1572 30528
rect 138 30408 1572 30442
rect 138 30322 1572 30356
rect 138 30236 1572 30270
rect 138 30150 1572 30184
rect 138 30064 1572 30098
rect 138 29978 1572 30012
rect 138 29892 1572 29926
rect 138 29806 1572 29840
rect 138 29720 1572 29754
rect 138 29634 1572 29668
rect 138 29548 1572 29582
rect 138 29462 1572 29496
rect 138 29376 1572 29410
rect 138 29290 1572 29324
rect 138 29204 1572 29238
rect 138 29118 1572 29152
rect 138 29032 1572 29066
rect 138 28946 1572 28980
rect 138 28860 1572 28894
rect 138 28774 1572 28808
rect 138 28688 1572 28722
rect 138 28602 1572 28636
rect 138 28516 1572 28550
rect 138 28430 1572 28464
rect 138 28344 1572 28378
rect 138 28258 1572 28292
rect 138 28172 1572 28206
rect 138 28086 1572 28120
rect 138 28000 1572 28034
rect 138 27914 1572 27948
rect 138 27828 1572 27862
rect 138 27742 1572 27776
rect 138 27656 1572 27690
rect 138 27570 1572 27604
rect 138 27484 1572 27518
rect 138 27398 1572 27432
rect 138 27312 1572 27346
rect 138 27226 1572 27260
rect 138 27140 1572 27174
rect 138 27054 1572 27088
rect 138 26968 1572 27002
rect 138 26882 1572 26916
rect 138 26796 1572 26830
rect 138 26710 1572 26744
rect 138 26624 1572 26658
rect 138 26538 1572 26572
rect 138 26452 1572 26486
rect 138 26366 1572 26400
rect 138 26280 1572 26314
rect 138 26194 1572 26228
rect 138 26108 1572 26142
rect 138 26022 1572 26056
rect 138 25936 1572 25970
rect 138 25850 1572 25884
rect 138 25764 1572 25798
rect 138 25678 1572 25712
rect 138 25592 1572 25626
rect 138 25506 1572 25540
rect 138 25420 1572 25454
rect 138 25334 1572 25368
rect 138 25248 1572 25282
rect 138 25162 1572 25196
rect 138 25076 1572 25110
rect 138 24990 1572 25024
rect 138 24904 1572 24938
rect 138 24818 1572 24852
rect 138 24732 1572 24766
rect 138 24646 1572 24680
rect 138 24560 1572 24594
rect 138 24474 1572 24508
rect 138 24388 1572 24422
rect 138 24302 1572 24336
rect 138 24216 1572 24250
rect 138 24130 1572 24164
rect 138 24044 1572 24078
rect 138 23958 1572 23992
rect 138 23872 1572 23906
rect 138 23786 1572 23820
rect 138 23700 1572 23734
rect 138 23614 1572 23648
rect 138 23528 1572 23562
rect 138 23442 1572 23476
rect 138 23356 1572 23390
rect 138 23270 1572 23304
rect 138 23184 1572 23218
rect 138 23098 1572 23132
rect 138 23012 1572 23046
rect 138 22926 1572 22960
rect 138 22840 1572 22874
rect 138 22754 1572 22788
rect 138 22668 1572 22702
rect 138 22582 1572 22616
rect 138 22496 1572 22530
rect 138 22410 1572 22444
rect 138 22324 1572 22358
rect 138 22238 1572 22272
rect 138 22152 1572 22186
rect 138 22066 1572 22100
rect 138 21980 1572 22014
rect 138 21894 1572 21928
rect 138 21808 1572 21842
rect 138 21722 1572 21756
rect 138 21636 1572 21670
rect 138 21550 1572 21584
rect 138 21464 1572 21498
rect 138 21378 1572 21412
rect 138 21292 1572 21326
rect 138 21206 1572 21240
rect 138 21120 1572 21154
rect 138 21034 1572 21068
rect 138 20948 1572 20982
rect 138 20862 1572 20896
rect 138 20776 1572 20810
rect 138 20690 1572 20724
rect 138 20604 1572 20638
rect 138 20518 1572 20552
rect 138 20432 1572 20466
rect 138 20346 1572 20380
rect 138 20260 1572 20294
rect 138 20174 1572 20208
rect 138 20088 1572 20122
rect 138 20002 1572 20036
rect 138 19916 1572 19950
rect 138 19830 1572 19864
rect 138 19744 1572 19778
rect 138 19658 1572 19692
rect 138 19572 1572 19606
rect 138 19486 1572 19520
rect 138 19400 1572 19434
rect 138 19314 1572 19348
rect 138 19228 1572 19262
rect 138 19142 1572 19176
rect 138 19056 1572 19090
rect 138 18970 1572 19004
rect 138 18884 1572 18918
rect 138 18798 1572 18832
rect 138 18712 1572 18746
rect 138 18626 1572 18660
rect 138 18540 1572 18574
rect 138 18454 1572 18488
rect 138 18368 1572 18402
rect 138 18282 1572 18316
rect 138 18196 1572 18230
rect 138 18110 1572 18144
rect 138 18024 1572 18058
rect 138 17938 1572 17972
rect 138 17852 1572 17886
rect 138 17766 1572 17800
rect 138 17680 1572 17714
rect 138 17594 1572 17628
rect 138 17508 1572 17542
rect 138 17422 1572 17456
rect 138 17336 1572 17370
rect 138 17250 1572 17284
rect 138 17164 1572 17198
rect 138 17078 1572 17112
rect 138 16992 1572 17026
rect 138 16906 1572 16940
rect 138 16820 1572 16854
rect 138 16734 1572 16768
rect 138 16648 1572 16682
rect 138 16562 1572 16596
rect 138 16476 1572 16510
rect 138 16390 1572 16424
rect 138 16304 1572 16338
rect 138 16218 1572 16252
rect 138 16132 1572 16166
rect 138 16046 1572 16080
rect 138 15960 1572 15994
rect 138 15874 1572 15908
rect 138 15788 1572 15822
rect 138 15702 1572 15736
rect 138 15616 1572 15650
rect 138 15530 1572 15564
rect 138 15444 1572 15478
rect 138 15358 1572 15392
rect 138 15272 1572 15306
rect 138 15186 1572 15220
rect 138 15100 1572 15134
rect 138 15014 1572 15048
rect 138 14928 1572 14962
rect 138 14842 1572 14876
rect 138 14756 1572 14790
rect 138 14670 1572 14704
rect 138 14584 1572 14618
rect 138 14498 1572 14532
rect 138 14412 1572 14446
rect 138 14326 1572 14360
rect 138 14240 1572 14274
rect 138 14154 1572 14188
rect 138 14068 1572 14102
rect 138 13982 1572 14016
rect 138 13896 1572 13930
rect 138 13810 1572 13844
rect 138 13724 1572 13758
rect 138 13638 1572 13672
rect 138 13552 1572 13586
rect 138 13466 1572 13500
rect 138 13380 1572 13414
rect 138 13294 1572 13328
rect 138 13208 1572 13242
rect 138 13122 1572 13156
rect 138 13036 1572 13070
rect 138 12950 1572 12984
rect 138 12864 1572 12898
rect 138 12778 1572 12812
rect 138 12692 1572 12726
rect 138 12606 1572 12640
rect 138 12520 1572 12554
rect 138 12434 1572 12468
rect 138 12348 1572 12382
rect 138 12262 1572 12296
rect 138 12176 1572 12210
rect 138 12090 1572 12124
rect 138 12004 1572 12038
rect 138 11918 1572 11952
rect 138 11832 1572 11866
rect 138 11746 1572 11780
rect 138 11660 1572 11694
rect 138 11574 1572 11608
rect 138 11488 1572 11522
rect 138 11402 1572 11436
rect 138 11316 1572 11350
rect 138 11230 1572 11264
rect 138 11144 1572 11178
rect 138 11058 1572 11092
rect 138 10972 1572 11006
rect 138 10886 1572 10920
rect 138 10800 1572 10834
rect 138 10714 1572 10748
rect 138 10628 1572 10662
rect 138 10542 1572 10576
rect 138 10456 1572 10490
rect 138 10370 1572 10404
rect 138 10284 1572 10318
rect 138 10198 1572 10232
rect 138 10112 1572 10146
rect 138 10026 1572 10060
rect 138 9940 1572 9974
rect 138 9854 1572 9888
rect 138 9768 1572 9802
rect 138 9682 1572 9716
rect 138 9596 1572 9630
rect 138 9510 1572 9544
rect 138 9424 1572 9458
rect 138 9338 1572 9372
rect 138 9252 1572 9286
rect 138 9166 1572 9200
rect 138 9080 1572 9114
rect 138 8994 1572 9028
rect 138 8908 1572 8942
rect 138 8822 1572 8856
rect 138 8736 1572 8770
rect 138 8650 1572 8684
rect 138 8564 1572 8598
rect 138 8478 1572 8512
rect 138 8392 1572 8426
rect 138 8306 1572 8340
rect 138 8220 1572 8254
rect 138 8134 1572 8168
rect 138 8048 1572 8082
rect 138 7962 1572 7996
rect 138 7876 1572 7910
rect 138 7790 1572 7824
rect 138 7704 1572 7738
rect 138 7618 1572 7652
rect 138 7532 1572 7566
rect 138 7446 1572 7480
rect 138 7360 1572 7394
rect 138 7274 1572 7308
rect 138 7188 1572 7222
rect 138 7102 1572 7136
rect 138 7016 1572 7050
rect 138 6930 1572 6964
rect 138 6844 1572 6878
rect 138 6758 1572 6792
rect 138 6672 1572 6706
rect 138 6586 1572 6620
rect 138 6500 1572 6534
rect 138 6414 1572 6448
rect 138 6328 1572 6362
rect 138 6242 1572 6276
rect 138 6156 1572 6190
rect 138 6070 1572 6104
rect 138 5984 1572 6018
rect 138 5898 1572 5932
rect 138 5812 1572 5846
rect 138 5726 1572 5760
rect 138 5640 1572 5674
rect 138 5554 1572 5588
rect 138 5468 1572 5502
rect 138 5382 1572 5416
rect 138 5296 1572 5330
rect 138 5210 1572 5244
rect 138 5124 1572 5158
rect 138 5038 1572 5072
rect 138 4952 1572 4986
rect 138 4866 1572 4900
rect 138 4780 1572 4814
rect 138 4694 1572 4728
rect 138 4608 1572 4642
rect 138 4522 1572 4556
rect 138 4436 1572 4470
rect 138 4350 1572 4384
rect 138 4264 1572 4298
rect 138 4178 1572 4212
rect 138 4092 1572 4126
rect 138 4006 1572 4040
rect 138 3920 1572 3954
rect 138 3834 1572 3868
rect 138 3748 1572 3782
rect 138 3662 1572 3696
rect 138 3576 1572 3610
rect 138 3490 1572 3524
rect 138 3404 1572 3438
rect 138 3318 1572 3352
rect 138 3232 1572 3266
rect 138 3146 1572 3180
rect 138 3060 1572 3094
rect 138 2974 1572 3008
rect 138 2888 1572 2922
rect 138 2802 1572 2836
rect 138 2716 1572 2750
rect 138 2630 1572 2664
rect 138 2544 1572 2578
rect 138 2458 1572 2492
rect 138 2372 1572 2406
rect 138 2286 1572 2320
rect 138 2200 1572 2234
rect 138 2114 1572 2148
rect 138 2028 1572 2062
rect 138 1942 1572 1976
rect 138 1856 1572 1890
rect 138 1770 1572 1804
rect 138 1684 1572 1718
rect 138 1598 1572 1632
rect 138 1512 1572 1546
rect 138 1426 1572 1460
rect 138 1340 1572 1374
rect 138 1254 1572 1288
rect 138 1168 1572 1202
rect 138 1082 1572 1116
rect 138 996 1572 1030
rect 138 910 1572 944
rect 138 824 1572 858
rect 138 738 1572 772
rect 138 652 1572 686
rect 138 566 1572 600
rect 138 480 1572 514
rect 138 394 1572 428
rect 138 308 1572 342
rect 138 222 1572 256
rect 1628 179 1662 43815
rect 138 136 1572 170
rect 1710 100 1744 43894
rect 100 36 1680 70
<< metal1 >>
rect 30 43958 1750 43964
rect 30 43924 100 43958
rect 1680 43924 1750 43958
rect 30 43918 1750 43924
rect 30 43894 76 43918
rect 30 100 36 43894
rect 70 100 76 43894
rect 1704 43894 1750 43918
rect 894 43864 900 43867
rect 126 43858 900 43864
rect 1548 43864 1554 43867
rect 1548 43858 1584 43864
rect 126 43824 138 43858
rect 1572 43824 1584 43858
rect 126 43818 900 43824
rect 894 43815 900 43818
rect 1548 43818 1584 43824
rect 1618 43825 1672 43831
rect 1548 43815 1554 43818
rect 156 43778 162 43781
rect 126 43772 162 43778
rect 810 43778 816 43781
rect 810 43772 1584 43778
rect 126 43738 138 43772
rect 1572 43738 1584 43772
rect 126 43732 162 43738
rect 156 43729 162 43732
rect 810 43732 1584 43738
rect 810 43729 816 43732
rect 894 43692 900 43695
rect 126 43686 900 43692
rect 1548 43692 1554 43695
rect 1548 43686 1584 43692
rect 126 43652 138 43686
rect 1572 43652 1584 43686
rect 126 43646 900 43652
rect 894 43643 900 43646
rect 1548 43646 1584 43652
rect 1548 43643 1554 43646
rect 156 43606 162 43609
rect 126 43600 162 43606
rect 810 43606 816 43609
rect 810 43600 1584 43606
rect 126 43566 138 43600
rect 1572 43566 1584 43600
rect 126 43560 162 43566
rect 156 43557 162 43560
rect 810 43560 1584 43566
rect 810 43557 816 43560
rect 894 43520 900 43523
rect 126 43514 900 43520
rect 1548 43520 1554 43523
rect 1548 43514 1584 43520
rect 126 43480 138 43514
rect 1572 43480 1584 43514
rect 126 43474 900 43480
rect 894 43471 900 43474
rect 1548 43474 1584 43480
rect 1548 43471 1554 43474
rect 156 43434 162 43437
rect 126 43428 162 43434
rect 810 43434 816 43437
rect 810 43428 1584 43434
rect 126 43394 138 43428
rect 1572 43394 1584 43428
rect 126 43388 162 43394
rect 156 43385 162 43388
rect 810 43388 1584 43394
rect 810 43385 816 43388
rect 894 43348 900 43351
rect 126 43342 900 43348
rect 1548 43348 1554 43351
rect 1548 43342 1584 43348
rect 126 43308 138 43342
rect 1572 43308 1584 43342
rect 126 43302 900 43308
rect 894 43299 900 43302
rect 1548 43302 1584 43308
rect 1548 43299 1554 43302
rect 156 43262 162 43265
rect 126 43256 162 43262
rect 810 43262 816 43265
rect 810 43256 1584 43262
rect 126 43222 138 43256
rect 1572 43222 1584 43256
rect 126 43216 162 43222
rect 156 43213 162 43216
rect 810 43216 1584 43222
rect 810 43213 816 43216
rect 894 43176 900 43179
rect 126 43170 900 43176
rect 1548 43176 1554 43179
rect 1548 43170 1584 43176
rect 126 43136 138 43170
rect 1572 43136 1584 43170
rect 126 43130 900 43136
rect 894 43127 900 43130
rect 1548 43130 1584 43136
rect 1548 43127 1554 43130
rect 156 43090 162 43093
rect 126 43084 162 43090
rect 810 43090 816 43093
rect 810 43084 1584 43090
rect 126 43050 138 43084
rect 1572 43050 1584 43084
rect 126 43044 162 43050
rect 156 43041 162 43044
rect 810 43044 1584 43050
rect 810 43041 816 43044
rect 894 43004 900 43007
rect 126 42998 900 43004
rect 1548 43004 1554 43007
rect 1548 42998 1584 43004
rect 126 42964 138 42998
rect 1572 42964 1584 42998
rect 126 42958 900 42964
rect 894 42955 900 42958
rect 1548 42958 1584 42964
rect 1548 42955 1554 42958
rect 156 42918 162 42921
rect 126 42912 162 42918
rect 810 42918 816 42921
rect 810 42912 1584 42918
rect 126 42878 138 42912
rect 1572 42878 1584 42912
rect 126 42872 162 42878
rect 156 42869 162 42872
rect 810 42872 1584 42878
rect 810 42869 816 42872
rect 894 42832 900 42835
rect 126 42826 900 42832
rect 1548 42832 1554 42835
rect 1548 42826 1584 42832
rect 126 42792 138 42826
rect 1572 42792 1584 42826
rect 126 42786 900 42792
rect 894 42783 900 42786
rect 1548 42786 1584 42792
rect 1548 42783 1554 42786
rect 156 42746 162 42749
rect 126 42740 162 42746
rect 810 42746 816 42749
rect 810 42740 1584 42746
rect 126 42706 138 42740
rect 1572 42706 1584 42740
rect 126 42700 162 42706
rect 156 42697 162 42700
rect 810 42700 1584 42706
rect 810 42697 816 42700
rect 894 42660 900 42663
rect 126 42654 900 42660
rect 1548 42660 1554 42663
rect 1548 42654 1584 42660
rect 126 42620 138 42654
rect 1572 42620 1584 42654
rect 126 42614 900 42620
rect 894 42611 900 42614
rect 1548 42614 1584 42620
rect 1548 42611 1554 42614
rect 156 42574 162 42577
rect 126 42568 162 42574
rect 810 42574 816 42577
rect 810 42568 1584 42574
rect 126 42534 138 42568
rect 1572 42534 1584 42568
rect 126 42528 162 42534
rect 156 42525 162 42528
rect 810 42528 1584 42534
rect 810 42525 816 42528
rect 894 42488 900 42491
rect 126 42482 900 42488
rect 1548 42488 1554 42491
rect 1548 42482 1584 42488
rect 126 42448 138 42482
rect 1572 42448 1584 42482
rect 126 42442 900 42448
rect 894 42439 900 42442
rect 1548 42442 1584 42448
rect 1548 42439 1554 42442
rect 156 42402 162 42405
rect 126 42396 162 42402
rect 810 42402 816 42405
rect 810 42396 1584 42402
rect 126 42362 138 42396
rect 1572 42362 1584 42396
rect 126 42356 162 42362
rect 156 42353 162 42356
rect 810 42356 1584 42362
rect 810 42353 816 42356
rect 894 42316 900 42319
rect 126 42310 900 42316
rect 1548 42316 1554 42319
rect 1548 42310 1584 42316
rect 126 42276 138 42310
rect 1572 42276 1584 42310
rect 126 42270 900 42276
rect 894 42267 900 42270
rect 1548 42270 1584 42276
rect 1548 42267 1554 42270
rect 156 42230 162 42233
rect 126 42224 162 42230
rect 810 42230 816 42233
rect 810 42224 1584 42230
rect 126 42190 138 42224
rect 1572 42190 1584 42224
rect 126 42184 162 42190
rect 156 42181 162 42184
rect 810 42184 1584 42190
rect 810 42181 816 42184
rect 894 42144 900 42147
rect 126 42138 900 42144
rect 1548 42144 1554 42147
rect 1548 42138 1584 42144
rect 126 42104 138 42138
rect 1572 42104 1584 42138
rect 126 42098 900 42104
rect 894 42095 900 42098
rect 1548 42098 1584 42104
rect 1548 42095 1554 42098
rect 156 42058 162 42061
rect 126 42052 162 42058
rect 810 42058 816 42061
rect 810 42052 1584 42058
rect 126 42018 138 42052
rect 1572 42018 1584 42052
rect 126 42012 162 42018
rect 156 42009 162 42012
rect 810 42012 1584 42018
rect 810 42009 816 42012
rect 894 41972 900 41975
rect 126 41966 900 41972
rect 1548 41972 1554 41975
rect 1548 41966 1584 41972
rect 126 41932 138 41966
rect 1572 41932 1584 41966
rect 126 41926 900 41932
rect 894 41923 900 41926
rect 1548 41926 1584 41932
rect 1548 41923 1554 41926
rect 156 41886 162 41889
rect 126 41880 162 41886
rect 810 41886 816 41889
rect 810 41880 1584 41886
rect 126 41846 138 41880
rect 1572 41846 1584 41880
rect 126 41840 162 41846
rect 156 41837 162 41840
rect 810 41840 1584 41846
rect 810 41837 816 41840
rect 894 41800 900 41803
rect 126 41794 900 41800
rect 1548 41800 1554 41803
rect 1548 41794 1584 41800
rect 126 41760 138 41794
rect 1572 41760 1584 41794
rect 126 41754 900 41760
rect 894 41751 900 41754
rect 1548 41754 1584 41760
rect 1548 41751 1554 41754
rect 156 41714 162 41717
rect 126 41708 162 41714
rect 810 41714 816 41717
rect 810 41708 1584 41714
rect 126 41674 138 41708
rect 1572 41674 1584 41708
rect 126 41668 162 41674
rect 156 41665 162 41668
rect 810 41668 1584 41674
rect 810 41665 816 41668
rect 894 41628 900 41631
rect 126 41622 900 41628
rect 1548 41628 1554 41631
rect 1548 41622 1584 41628
rect 126 41588 138 41622
rect 1572 41588 1584 41622
rect 126 41582 900 41588
rect 894 41579 900 41582
rect 1548 41582 1584 41588
rect 1548 41579 1554 41582
rect 156 41542 162 41545
rect 126 41536 162 41542
rect 810 41542 816 41545
rect 810 41536 1584 41542
rect 126 41502 138 41536
rect 1572 41502 1584 41536
rect 126 41496 162 41502
rect 156 41493 162 41496
rect 810 41496 1584 41502
rect 810 41493 816 41496
rect 894 41456 900 41459
rect 126 41450 900 41456
rect 1548 41456 1554 41459
rect 1548 41450 1584 41456
rect 126 41416 138 41450
rect 1572 41416 1584 41450
rect 126 41410 900 41416
rect 894 41407 900 41410
rect 1548 41410 1584 41416
rect 1548 41407 1554 41410
rect 156 41370 162 41373
rect 126 41364 162 41370
rect 810 41370 816 41373
rect 810 41364 1584 41370
rect 126 41330 138 41364
rect 1572 41330 1584 41364
rect 126 41324 162 41330
rect 156 41321 162 41324
rect 810 41324 1584 41330
rect 810 41321 816 41324
rect 894 41284 900 41287
rect 126 41278 900 41284
rect 1548 41284 1554 41287
rect 1548 41278 1584 41284
rect 126 41244 138 41278
rect 1572 41244 1584 41278
rect 126 41238 900 41244
rect 894 41235 900 41238
rect 1548 41238 1584 41244
rect 1548 41235 1554 41238
rect 156 41198 162 41201
rect 126 41192 162 41198
rect 810 41198 816 41201
rect 810 41192 1584 41198
rect 126 41158 138 41192
rect 1572 41158 1584 41192
rect 126 41152 162 41158
rect 156 41149 162 41152
rect 810 41152 1584 41158
rect 810 41149 816 41152
rect 894 41112 900 41115
rect 126 41106 900 41112
rect 1548 41112 1554 41115
rect 1548 41106 1584 41112
rect 126 41072 138 41106
rect 1572 41072 1584 41106
rect 126 41066 900 41072
rect 894 41063 900 41066
rect 1548 41066 1584 41072
rect 1548 41063 1554 41066
rect 156 41026 162 41029
rect 126 41020 162 41026
rect 810 41026 816 41029
rect 810 41020 1584 41026
rect 126 40986 138 41020
rect 1572 40986 1584 41020
rect 126 40980 162 40986
rect 156 40977 162 40980
rect 810 40980 1584 40986
rect 810 40977 816 40980
rect 894 40940 900 40943
rect 126 40934 900 40940
rect 1548 40940 1554 40943
rect 1548 40934 1584 40940
rect 126 40900 138 40934
rect 1572 40900 1584 40934
rect 126 40894 900 40900
rect 894 40891 900 40894
rect 1548 40894 1584 40900
rect 1548 40891 1554 40894
rect 156 40854 162 40857
rect 126 40848 162 40854
rect 810 40854 816 40857
rect 810 40848 1584 40854
rect 126 40814 138 40848
rect 1572 40814 1584 40848
rect 126 40808 162 40814
rect 156 40805 162 40808
rect 810 40808 1584 40814
rect 810 40805 816 40808
rect 894 40768 900 40771
rect 126 40762 900 40768
rect 1548 40768 1554 40771
rect 1548 40762 1584 40768
rect 126 40728 138 40762
rect 1572 40728 1584 40762
rect 126 40722 900 40728
rect 894 40719 900 40722
rect 1548 40722 1584 40728
rect 1548 40719 1554 40722
rect 156 40682 162 40685
rect 126 40676 162 40682
rect 810 40682 816 40685
rect 810 40676 1584 40682
rect 126 40642 138 40676
rect 1572 40642 1584 40676
rect 126 40636 162 40642
rect 156 40633 162 40636
rect 810 40636 1584 40642
rect 810 40633 816 40636
rect 894 40596 900 40599
rect 126 40590 900 40596
rect 1548 40596 1554 40599
rect 1548 40590 1584 40596
rect 126 40556 138 40590
rect 1572 40556 1584 40590
rect 126 40550 900 40556
rect 894 40547 900 40550
rect 1548 40550 1584 40556
rect 1548 40547 1554 40550
rect 156 40510 162 40513
rect 126 40504 162 40510
rect 810 40510 816 40513
rect 810 40504 1584 40510
rect 126 40470 138 40504
rect 1572 40470 1584 40504
rect 126 40464 162 40470
rect 156 40461 162 40464
rect 810 40464 1584 40470
rect 810 40461 816 40464
rect 894 40424 900 40427
rect 126 40418 900 40424
rect 1548 40424 1554 40427
rect 1548 40418 1584 40424
rect 126 40384 138 40418
rect 1572 40384 1584 40418
rect 126 40378 900 40384
rect 894 40375 900 40378
rect 1548 40378 1584 40384
rect 1548 40375 1554 40378
rect 156 40338 162 40341
rect 126 40332 162 40338
rect 810 40338 816 40341
rect 810 40332 1584 40338
rect 126 40298 138 40332
rect 1572 40298 1584 40332
rect 126 40292 162 40298
rect 156 40289 162 40292
rect 810 40292 1584 40298
rect 810 40289 816 40292
rect 894 40252 900 40255
rect 126 40246 900 40252
rect 1548 40252 1554 40255
rect 1548 40246 1584 40252
rect 126 40212 138 40246
rect 1572 40212 1584 40246
rect 126 40206 900 40212
rect 894 40203 900 40206
rect 1548 40206 1584 40212
rect 1548 40203 1554 40206
rect 156 40166 162 40169
rect 126 40160 162 40166
rect 810 40166 816 40169
rect 810 40160 1584 40166
rect 126 40126 138 40160
rect 1572 40126 1584 40160
rect 126 40120 162 40126
rect 156 40117 162 40120
rect 810 40120 1584 40126
rect 810 40117 816 40120
rect 894 40080 900 40083
rect 126 40074 900 40080
rect 1548 40080 1554 40083
rect 1548 40074 1584 40080
rect 126 40040 138 40074
rect 1572 40040 1584 40074
rect 126 40034 900 40040
rect 894 40031 900 40034
rect 1548 40034 1584 40040
rect 1548 40031 1554 40034
rect 156 39994 162 39997
rect 126 39988 162 39994
rect 810 39994 816 39997
rect 810 39988 1584 39994
rect 126 39954 138 39988
rect 1572 39954 1584 39988
rect 126 39948 162 39954
rect 156 39945 162 39948
rect 810 39948 1584 39954
rect 810 39945 816 39948
rect 894 39908 900 39911
rect 126 39902 900 39908
rect 1548 39908 1554 39911
rect 1548 39902 1584 39908
rect 126 39868 138 39902
rect 1572 39868 1584 39902
rect 126 39862 900 39868
rect 894 39859 900 39862
rect 1548 39862 1584 39868
rect 1548 39859 1554 39862
rect 156 39822 162 39825
rect 126 39816 162 39822
rect 810 39822 816 39825
rect 810 39816 1584 39822
rect 126 39782 138 39816
rect 1572 39782 1584 39816
rect 126 39776 162 39782
rect 156 39773 162 39776
rect 810 39776 1584 39782
rect 810 39773 816 39776
rect 894 39736 900 39739
rect 126 39730 900 39736
rect 1548 39736 1554 39739
rect 1548 39730 1584 39736
rect 126 39696 138 39730
rect 1572 39696 1584 39730
rect 126 39690 900 39696
rect 894 39687 900 39690
rect 1548 39690 1584 39696
rect 1548 39687 1554 39690
rect 156 39650 162 39653
rect 126 39644 162 39650
rect 810 39650 816 39653
rect 810 39644 1584 39650
rect 126 39610 138 39644
rect 1572 39610 1584 39644
rect 126 39604 162 39610
rect 156 39601 162 39604
rect 810 39604 1584 39610
rect 810 39601 816 39604
rect 894 39564 900 39567
rect 126 39558 900 39564
rect 1548 39564 1554 39567
rect 1548 39558 1584 39564
rect 126 39524 138 39558
rect 1572 39524 1584 39558
rect 126 39518 900 39524
rect 894 39515 900 39518
rect 1548 39518 1584 39524
rect 1548 39515 1554 39518
rect 156 39478 162 39481
rect 126 39472 162 39478
rect 810 39478 816 39481
rect 810 39472 1584 39478
rect 126 39438 138 39472
rect 1572 39438 1584 39472
rect 126 39432 162 39438
rect 156 39429 162 39432
rect 810 39432 1584 39438
rect 810 39429 816 39432
rect 894 39392 900 39395
rect 126 39386 900 39392
rect 1548 39392 1554 39395
rect 1548 39386 1584 39392
rect 126 39352 138 39386
rect 1572 39352 1584 39386
rect 126 39346 900 39352
rect 894 39343 900 39346
rect 1548 39346 1584 39352
rect 1548 39343 1554 39346
rect 156 39306 162 39309
rect 126 39300 162 39306
rect 810 39306 816 39309
rect 810 39300 1584 39306
rect 126 39266 138 39300
rect 1572 39266 1584 39300
rect 126 39260 162 39266
rect 156 39257 162 39260
rect 810 39260 1584 39266
rect 810 39257 816 39260
rect 894 39220 900 39223
rect 126 39214 900 39220
rect 1548 39220 1554 39223
rect 1548 39214 1584 39220
rect 126 39180 138 39214
rect 1572 39180 1584 39214
rect 126 39174 900 39180
rect 894 39171 900 39174
rect 1548 39174 1584 39180
rect 1548 39171 1554 39174
rect 156 39134 162 39137
rect 126 39128 162 39134
rect 810 39134 816 39137
rect 810 39128 1584 39134
rect 126 39094 138 39128
rect 1572 39094 1584 39128
rect 126 39088 162 39094
rect 156 39085 162 39088
rect 810 39088 1584 39094
rect 810 39085 816 39088
rect 894 39048 900 39051
rect 126 39042 900 39048
rect 1548 39048 1554 39051
rect 1548 39042 1584 39048
rect 126 39008 138 39042
rect 1572 39008 1584 39042
rect 126 39002 900 39008
rect 894 38999 900 39002
rect 1548 39002 1584 39008
rect 1548 38999 1554 39002
rect 156 38962 162 38965
rect 126 38956 162 38962
rect 810 38962 816 38965
rect 810 38956 1584 38962
rect 126 38922 138 38956
rect 1572 38922 1584 38956
rect 126 38916 162 38922
rect 156 38913 162 38916
rect 810 38916 1584 38922
rect 810 38913 816 38916
rect 894 38876 900 38879
rect 126 38870 900 38876
rect 1548 38876 1554 38879
rect 1548 38870 1584 38876
rect 126 38836 138 38870
rect 1572 38836 1584 38870
rect 126 38830 900 38836
rect 894 38827 900 38830
rect 1548 38830 1584 38836
rect 1548 38827 1554 38830
rect 156 38790 162 38793
rect 126 38784 162 38790
rect 810 38790 816 38793
rect 810 38784 1584 38790
rect 126 38750 138 38784
rect 1572 38750 1584 38784
rect 126 38744 162 38750
rect 156 38741 162 38744
rect 810 38744 1584 38750
rect 810 38741 816 38744
rect 894 38704 900 38707
rect 126 38698 900 38704
rect 1548 38704 1554 38707
rect 1548 38698 1584 38704
rect 126 38664 138 38698
rect 1572 38664 1584 38698
rect 126 38658 900 38664
rect 894 38655 900 38658
rect 1548 38658 1584 38664
rect 1548 38655 1554 38658
rect 156 38618 162 38621
rect 126 38612 162 38618
rect 810 38618 816 38621
rect 810 38612 1584 38618
rect 126 38578 138 38612
rect 1572 38578 1584 38612
rect 126 38572 162 38578
rect 156 38569 162 38572
rect 810 38572 1584 38578
rect 810 38569 816 38572
rect 894 38532 900 38535
rect 126 38526 900 38532
rect 1548 38532 1554 38535
rect 1548 38526 1584 38532
rect 126 38492 138 38526
rect 1572 38492 1584 38526
rect 126 38486 900 38492
rect 894 38483 900 38486
rect 1548 38486 1584 38492
rect 1548 38483 1554 38486
rect 156 38446 162 38449
rect 126 38440 162 38446
rect 810 38446 816 38449
rect 810 38440 1584 38446
rect 126 38406 138 38440
rect 1572 38406 1584 38440
rect 126 38400 162 38406
rect 156 38397 162 38400
rect 810 38400 1584 38406
rect 810 38397 816 38400
rect 894 38360 900 38363
rect 126 38354 900 38360
rect 1548 38360 1554 38363
rect 1548 38354 1584 38360
rect 126 38320 138 38354
rect 1572 38320 1584 38354
rect 126 38314 900 38320
rect 894 38311 900 38314
rect 1548 38314 1584 38320
rect 1548 38311 1554 38314
rect 156 38274 162 38277
rect 126 38268 162 38274
rect 810 38274 816 38277
rect 810 38268 1584 38274
rect 126 38234 138 38268
rect 1572 38234 1584 38268
rect 126 38228 162 38234
rect 156 38225 162 38228
rect 810 38228 1584 38234
rect 810 38225 816 38228
rect 894 38188 900 38191
rect 126 38182 900 38188
rect 1548 38188 1554 38191
rect 1548 38182 1584 38188
rect 126 38148 138 38182
rect 1572 38148 1584 38182
rect 126 38142 900 38148
rect 894 38139 900 38142
rect 1548 38142 1584 38148
rect 1548 38139 1554 38142
rect 156 38102 162 38105
rect 126 38096 162 38102
rect 810 38102 816 38105
rect 810 38096 1584 38102
rect 126 38062 138 38096
rect 1572 38062 1584 38096
rect 126 38056 162 38062
rect 156 38053 162 38056
rect 810 38056 1584 38062
rect 810 38053 816 38056
rect 894 38016 900 38019
rect 126 38010 900 38016
rect 1548 38016 1554 38019
rect 1548 38010 1584 38016
rect 126 37976 138 38010
rect 1572 37976 1584 38010
rect 126 37970 900 37976
rect 894 37967 900 37970
rect 1548 37970 1584 37976
rect 1548 37967 1554 37970
rect 156 37930 162 37933
rect 126 37924 162 37930
rect 810 37930 816 37933
rect 810 37924 1584 37930
rect 126 37890 138 37924
rect 1572 37890 1584 37924
rect 126 37884 162 37890
rect 156 37881 162 37884
rect 810 37884 1584 37890
rect 810 37881 816 37884
rect 894 37844 900 37847
rect 126 37838 900 37844
rect 1548 37844 1554 37847
rect 1548 37838 1584 37844
rect 126 37804 138 37838
rect 1572 37804 1584 37838
rect 126 37798 900 37804
rect 894 37795 900 37798
rect 1548 37798 1584 37804
rect 1548 37795 1554 37798
rect 156 37758 162 37761
rect 126 37752 162 37758
rect 810 37758 816 37761
rect 810 37752 1584 37758
rect 126 37718 138 37752
rect 1572 37718 1584 37752
rect 126 37712 162 37718
rect 156 37709 162 37712
rect 810 37712 1584 37718
rect 810 37709 816 37712
rect 894 37672 900 37675
rect 126 37666 900 37672
rect 1548 37672 1554 37675
rect 1548 37666 1584 37672
rect 126 37632 138 37666
rect 1572 37632 1584 37666
rect 126 37626 900 37632
rect 894 37623 900 37626
rect 1548 37626 1584 37632
rect 1548 37623 1554 37626
rect 156 37586 162 37589
rect 126 37580 162 37586
rect 810 37586 816 37589
rect 810 37580 1584 37586
rect 126 37546 138 37580
rect 1572 37546 1584 37580
rect 126 37540 162 37546
rect 156 37537 162 37540
rect 810 37540 1584 37546
rect 810 37537 816 37540
rect 894 37500 900 37503
rect 126 37494 900 37500
rect 1548 37500 1554 37503
rect 1548 37494 1584 37500
rect 126 37460 138 37494
rect 1572 37460 1584 37494
rect 126 37454 900 37460
rect 894 37451 900 37454
rect 1548 37454 1584 37460
rect 1548 37451 1554 37454
rect 156 37414 162 37417
rect 126 37408 162 37414
rect 810 37414 816 37417
rect 810 37408 1584 37414
rect 126 37374 138 37408
rect 1572 37374 1584 37408
rect 126 37368 162 37374
rect 156 37365 162 37368
rect 810 37368 1584 37374
rect 810 37365 816 37368
rect 894 37328 900 37331
rect 126 37322 900 37328
rect 1548 37328 1554 37331
rect 1548 37322 1584 37328
rect 126 37288 138 37322
rect 1572 37288 1584 37322
rect 126 37282 900 37288
rect 894 37279 900 37282
rect 1548 37282 1584 37288
rect 1548 37279 1554 37282
rect 156 37242 162 37245
rect 126 37236 162 37242
rect 810 37242 816 37245
rect 810 37236 1584 37242
rect 126 37202 138 37236
rect 1572 37202 1584 37236
rect 126 37196 162 37202
rect 156 37193 162 37196
rect 810 37196 1584 37202
rect 810 37193 816 37196
rect 894 37156 900 37159
rect 126 37150 900 37156
rect 1548 37156 1554 37159
rect 1548 37150 1584 37156
rect 126 37116 138 37150
rect 1572 37116 1584 37150
rect 126 37110 900 37116
rect 894 37107 900 37110
rect 1548 37110 1584 37116
rect 1548 37107 1554 37110
rect 156 37070 162 37073
rect 126 37064 162 37070
rect 810 37070 816 37073
rect 810 37064 1584 37070
rect 126 37030 138 37064
rect 1572 37030 1584 37064
rect 126 37024 162 37030
rect 156 37021 162 37024
rect 810 37024 1584 37030
rect 810 37021 816 37024
rect 894 36984 900 36987
rect 126 36978 900 36984
rect 1548 36984 1554 36987
rect 1548 36978 1584 36984
rect 126 36944 138 36978
rect 1572 36944 1584 36978
rect 126 36938 900 36944
rect 894 36935 900 36938
rect 1548 36938 1584 36944
rect 1548 36935 1554 36938
rect 156 36898 162 36901
rect 126 36892 162 36898
rect 810 36898 816 36901
rect 810 36892 1584 36898
rect 126 36858 138 36892
rect 1572 36858 1584 36892
rect 126 36852 162 36858
rect 156 36849 162 36852
rect 810 36852 1584 36858
rect 810 36849 816 36852
rect 894 36812 900 36815
rect 126 36806 900 36812
rect 1548 36812 1554 36815
rect 1548 36806 1584 36812
rect 126 36772 138 36806
rect 1572 36772 1584 36806
rect 126 36766 900 36772
rect 894 36763 900 36766
rect 1548 36766 1584 36772
rect 1548 36763 1554 36766
rect 156 36726 162 36729
rect 126 36720 162 36726
rect 810 36726 816 36729
rect 810 36720 1584 36726
rect 126 36686 138 36720
rect 1572 36686 1584 36720
rect 126 36680 162 36686
rect 156 36677 162 36680
rect 810 36680 1584 36686
rect 810 36677 816 36680
rect 894 36640 900 36643
rect 126 36634 900 36640
rect 1548 36640 1554 36643
rect 1548 36634 1584 36640
rect 126 36600 138 36634
rect 1572 36600 1584 36634
rect 126 36594 900 36600
rect 894 36591 900 36594
rect 1548 36594 1584 36600
rect 1548 36591 1554 36594
rect 156 36554 162 36557
rect 126 36548 162 36554
rect 810 36554 816 36557
rect 810 36548 1584 36554
rect 126 36514 138 36548
rect 1572 36514 1584 36548
rect 126 36508 162 36514
rect 156 36505 162 36508
rect 810 36508 1584 36514
rect 810 36505 816 36508
rect 894 36468 900 36471
rect 126 36462 900 36468
rect 1548 36468 1554 36471
rect 1548 36462 1584 36468
rect 126 36428 138 36462
rect 1572 36428 1584 36462
rect 126 36422 900 36428
rect 894 36419 900 36422
rect 1548 36422 1584 36428
rect 1548 36419 1554 36422
rect 156 36382 162 36385
rect 126 36376 162 36382
rect 810 36382 816 36385
rect 810 36376 1584 36382
rect 126 36342 138 36376
rect 1572 36342 1584 36376
rect 126 36336 162 36342
rect 156 36333 162 36336
rect 810 36336 1584 36342
rect 810 36333 816 36336
rect 894 36296 900 36299
rect 126 36290 900 36296
rect 1548 36296 1554 36299
rect 1548 36290 1584 36296
rect 126 36256 138 36290
rect 1572 36256 1584 36290
rect 126 36250 900 36256
rect 894 36247 900 36250
rect 1548 36250 1584 36256
rect 1548 36247 1554 36250
rect 156 36210 162 36213
rect 126 36204 162 36210
rect 810 36210 816 36213
rect 810 36204 1584 36210
rect 126 36170 138 36204
rect 1572 36170 1584 36204
rect 126 36164 162 36170
rect 156 36161 162 36164
rect 810 36164 1584 36170
rect 810 36161 816 36164
rect 894 36124 900 36127
rect 126 36118 900 36124
rect 1548 36124 1554 36127
rect 1548 36118 1584 36124
rect 126 36084 138 36118
rect 1572 36084 1584 36118
rect 126 36078 900 36084
rect 894 36075 900 36078
rect 1548 36078 1584 36084
rect 1548 36075 1554 36078
rect 156 36038 162 36041
rect 126 36032 162 36038
rect 810 36038 816 36041
rect 810 36032 1584 36038
rect 126 35998 138 36032
rect 1572 35998 1584 36032
rect 126 35992 162 35998
rect 156 35989 162 35992
rect 810 35992 1584 35998
rect 810 35989 816 35992
rect 894 35952 900 35955
rect 126 35946 900 35952
rect 1548 35952 1554 35955
rect 1548 35946 1584 35952
rect 126 35912 138 35946
rect 1572 35912 1584 35946
rect 126 35906 900 35912
rect 894 35903 900 35906
rect 1548 35906 1584 35912
rect 1548 35903 1554 35906
rect 156 35866 162 35869
rect 126 35860 162 35866
rect 810 35866 816 35869
rect 810 35860 1584 35866
rect 126 35826 138 35860
rect 1572 35826 1584 35860
rect 126 35820 162 35826
rect 156 35817 162 35820
rect 810 35820 1584 35826
rect 810 35817 816 35820
rect 894 35780 900 35783
rect 126 35774 900 35780
rect 1548 35780 1554 35783
rect 1548 35774 1584 35780
rect 126 35740 138 35774
rect 1572 35740 1584 35774
rect 126 35734 900 35740
rect 894 35731 900 35734
rect 1548 35734 1584 35740
rect 1548 35731 1554 35734
rect 156 35694 162 35697
rect 126 35688 162 35694
rect 810 35694 816 35697
rect 810 35688 1584 35694
rect 126 35654 138 35688
rect 1572 35654 1584 35688
rect 126 35648 162 35654
rect 156 35645 162 35648
rect 810 35648 1584 35654
rect 810 35645 816 35648
rect 894 35608 900 35611
rect 126 35602 900 35608
rect 1548 35608 1554 35611
rect 1548 35602 1584 35608
rect 126 35568 138 35602
rect 1572 35568 1584 35602
rect 126 35562 900 35568
rect 894 35559 900 35562
rect 1548 35562 1584 35568
rect 1548 35559 1554 35562
rect 156 35522 162 35525
rect 126 35516 162 35522
rect 810 35522 816 35525
rect 810 35516 1584 35522
rect 126 35482 138 35516
rect 1572 35482 1584 35516
rect 126 35476 162 35482
rect 156 35473 162 35476
rect 810 35476 1584 35482
rect 810 35473 816 35476
rect 894 35436 900 35439
rect 126 35430 900 35436
rect 1548 35436 1554 35439
rect 1548 35430 1584 35436
rect 126 35396 138 35430
rect 1572 35396 1584 35430
rect 126 35390 900 35396
rect 894 35387 900 35390
rect 1548 35390 1584 35396
rect 1548 35387 1554 35390
rect 156 35350 162 35353
rect 126 35344 162 35350
rect 810 35350 816 35353
rect 810 35344 1584 35350
rect 126 35310 138 35344
rect 1572 35310 1584 35344
rect 126 35304 162 35310
rect 156 35301 162 35304
rect 810 35304 1584 35310
rect 810 35301 816 35304
rect 894 35264 900 35267
rect 126 35258 900 35264
rect 1548 35264 1554 35267
rect 1548 35258 1584 35264
rect 126 35224 138 35258
rect 1572 35224 1584 35258
rect 126 35218 900 35224
rect 894 35215 900 35218
rect 1548 35218 1584 35224
rect 1548 35215 1554 35218
rect 156 35178 162 35181
rect 126 35172 162 35178
rect 810 35178 816 35181
rect 810 35172 1584 35178
rect 126 35138 138 35172
rect 1572 35138 1584 35172
rect 126 35132 162 35138
rect 156 35129 162 35132
rect 810 35132 1584 35138
rect 810 35129 816 35132
rect 894 35092 900 35095
rect 126 35086 900 35092
rect 1548 35092 1554 35095
rect 1548 35086 1584 35092
rect 126 35052 138 35086
rect 1572 35052 1584 35086
rect 126 35046 900 35052
rect 894 35043 900 35046
rect 1548 35046 1584 35052
rect 1548 35043 1554 35046
rect 156 35006 162 35009
rect 126 35000 162 35006
rect 810 35006 816 35009
rect 810 35000 1584 35006
rect 126 34966 138 35000
rect 1572 34966 1584 35000
rect 126 34960 162 34966
rect 156 34957 162 34960
rect 810 34960 1584 34966
rect 810 34957 816 34960
rect 894 34920 900 34923
rect 126 34914 900 34920
rect 1548 34920 1554 34923
rect 1548 34914 1584 34920
rect 126 34880 138 34914
rect 1572 34880 1584 34914
rect 126 34874 900 34880
rect 894 34871 900 34874
rect 1548 34874 1584 34880
rect 1548 34871 1554 34874
rect 156 34834 162 34837
rect 126 34828 162 34834
rect 810 34834 816 34837
rect 810 34828 1584 34834
rect 126 34794 138 34828
rect 1572 34794 1584 34828
rect 126 34788 162 34794
rect 156 34785 162 34788
rect 810 34788 1584 34794
rect 810 34785 816 34788
rect 894 34748 900 34751
rect 126 34742 900 34748
rect 1548 34748 1554 34751
rect 1548 34742 1584 34748
rect 126 34708 138 34742
rect 1572 34708 1584 34742
rect 126 34702 900 34708
rect 894 34699 900 34702
rect 1548 34702 1584 34708
rect 1548 34699 1554 34702
rect 156 34662 162 34665
rect 126 34656 162 34662
rect 810 34662 816 34665
rect 810 34656 1584 34662
rect 126 34622 138 34656
rect 1572 34622 1584 34656
rect 126 34616 162 34622
rect 156 34613 162 34616
rect 810 34616 1584 34622
rect 810 34613 816 34616
rect 894 34576 900 34579
rect 126 34570 900 34576
rect 1548 34576 1554 34579
rect 1548 34570 1584 34576
rect 126 34536 138 34570
rect 1572 34536 1584 34570
rect 126 34530 900 34536
rect 894 34527 900 34530
rect 1548 34530 1584 34536
rect 1548 34527 1554 34530
rect 156 34490 162 34493
rect 126 34484 162 34490
rect 810 34490 816 34493
rect 810 34484 1584 34490
rect 126 34450 138 34484
rect 1572 34450 1584 34484
rect 126 34444 162 34450
rect 156 34441 162 34444
rect 810 34444 1584 34450
rect 810 34441 816 34444
rect 894 34404 900 34407
rect 126 34398 900 34404
rect 1548 34404 1554 34407
rect 1548 34398 1584 34404
rect 126 34364 138 34398
rect 1572 34364 1584 34398
rect 126 34358 900 34364
rect 894 34355 900 34358
rect 1548 34358 1584 34364
rect 1548 34355 1554 34358
rect 156 34318 162 34321
rect 126 34312 162 34318
rect 810 34318 816 34321
rect 810 34312 1584 34318
rect 126 34278 138 34312
rect 1572 34278 1584 34312
rect 126 34272 162 34278
rect 156 34269 162 34272
rect 810 34272 1584 34278
rect 810 34269 816 34272
rect 894 34232 900 34235
rect 126 34226 900 34232
rect 1548 34232 1554 34235
rect 1548 34226 1584 34232
rect 126 34192 138 34226
rect 1572 34192 1584 34226
rect 126 34186 900 34192
rect 894 34183 900 34186
rect 1548 34186 1584 34192
rect 1548 34183 1554 34186
rect 156 34146 162 34149
rect 126 34140 162 34146
rect 810 34146 816 34149
rect 810 34140 1584 34146
rect 126 34106 138 34140
rect 1572 34106 1584 34140
rect 126 34100 162 34106
rect 156 34097 162 34100
rect 810 34100 1584 34106
rect 810 34097 816 34100
rect 894 34060 900 34063
rect 126 34054 900 34060
rect 1548 34060 1554 34063
rect 1548 34054 1584 34060
rect 126 34020 138 34054
rect 1572 34020 1584 34054
rect 126 34014 900 34020
rect 894 34011 900 34014
rect 1548 34014 1584 34020
rect 1548 34011 1554 34014
rect 156 33974 162 33977
rect 126 33968 162 33974
rect 810 33974 816 33977
rect 810 33968 1584 33974
rect 126 33934 138 33968
rect 1572 33934 1584 33968
rect 126 33928 162 33934
rect 156 33925 162 33928
rect 810 33928 1584 33934
rect 810 33925 816 33928
rect 894 33888 900 33891
rect 126 33882 900 33888
rect 1548 33888 1554 33891
rect 1548 33882 1584 33888
rect 126 33848 138 33882
rect 1572 33848 1584 33882
rect 126 33842 900 33848
rect 894 33839 900 33842
rect 1548 33842 1584 33848
rect 1548 33839 1554 33842
rect 156 33802 162 33805
rect 126 33796 162 33802
rect 810 33802 816 33805
rect 810 33796 1584 33802
rect 126 33762 138 33796
rect 1572 33762 1584 33796
rect 126 33756 162 33762
rect 156 33753 162 33756
rect 810 33756 1584 33762
rect 810 33753 816 33756
rect 894 33716 900 33719
rect 126 33710 900 33716
rect 1548 33716 1554 33719
rect 1548 33710 1584 33716
rect 126 33676 138 33710
rect 1572 33676 1584 33710
rect 126 33670 900 33676
rect 894 33667 900 33670
rect 1548 33670 1584 33676
rect 1548 33667 1554 33670
rect 156 33630 162 33633
rect 126 33624 162 33630
rect 810 33630 816 33633
rect 810 33624 1584 33630
rect 126 33590 138 33624
rect 1572 33590 1584 33624
rect 126 33584 162 33590
rect 156 33581 162 33584
rect 810 33584 1584 33590
rect 810 33581 816 33584
rect 894 33544 900 33547
rect 126 33538 900 33544
rect 1548 33544 1554 33547
rect 1548 33538 1584 33544
rect 126 33504 138 33538
rect 1572 33504 1584 33538
rect 126 33498 900 33504
rect 894 33495 900 33498
rect 1548 33498 1584 33504
rect 1548 33495 1554 33498
rect 156 33458 162 33461
rect 126 33452 162 33458
rect 810 33458 816 33461
rect 810 33452 1584 33458
rect 126 33418 138 33452
rect 1572 33418 1584 33452
rect 126 33412 162 33418
rect 156 33409 162 33412
rect 810 33412 1584 33418
rect 810 33409 816 33412
rect 894 33372 900 33375
rect 126 33366 900 33372
rect 1548 33372 1554 33375
rect 1548 33366 1584 33372
rect 126 33332 138 33366
rect 1572 33332 1584 33366
rect 126 33326 900 33332
rect 894 33323 900 33326
rect 1548 33326 1584 33332
rect 1548 33323 1554 33326
rect 156 33286 162 33289
rect 126 33280 162 33286
rect 810 33286 816 33289
rect 810 33280 1584 33286
rect 126 33246 138 33280
rect 1572 33246 1584 33280
rect 126 33240 162 33246
rect 156 33237 162 33240
rect 810 33240 1584 33246
rect 810 33237 816 33240
rect 894 33200 900 33203
rect 126 33194 900 33200
rect 1548 33200 1554 33203
rect 1548 33194 1584 33200
rect 126 33160 138 33194
rect 1572 33160 1584 33194
rect 126 33154 900 33160
rect 894 33151 900 33154
rect 1548 33154 1584 33160
rect 1548 33151 1554 33154
rect 156 33114 162 33117
rect 126 33108 162 33114
rect 810 33114 816 33117
rect 810 33108 1584 33114
rect 126 33074 138 33108
rect 1572 33074 1584 33108
rect 126 33068 162 33074
rect 156 33065 162 33068
rect 810 33068 1584 33074
rect 810 33065 816 33068
rect 894 33028 900 33031
rect 126 33022 900 33028
rect 1548 33028 1554 33031
rect 1548 33022 1584 33028
rect 126 32988 138 33022
rect 1572 32988 1584 33022
rect 126 32982 900 32988
rect 894 32979 900 32982
rect 1548 32982 1584 32988
rect 1548 32979 1554 32982
rect 156 32942 162 32945
rect 126 32936 162 32942
rect 810 32942 816 32945
rect 810 32936 1584 32942
rect 126 32902 138 32936
rect 1572 32902 1584 32936
rect 126 32896 162 32902
rect 156 32893 162 32896
rect 810 32896 1584 32902
rect 810 32893 816 32896
rect 894 32856 900 32859
rect 126 32850 900 32856
rect 1548 32856 1554 32859
rect 1548 32850 1584 32856
rect 126 32816 138 32850
rect 1572 32816 1584 32850
rect 126 32810 900 32816
rect 894 32807 900 32810
rect 1548 32810 1584 32816
rect 1548 32807 1554 32810
rect 156 32770 162 32773
rect 126 32764 162 32770
rect 810 32770 816 32773
rect 810 32764 1584 32770
rect 126 32730 138 32764
rect 1572 32730 1584 32764
rect 126 32724 162 32730
rect 156 32721 162 32724
rect 810 32724 1584 32730
rect 810 32721 816 32724
rect 894 32684 900 32687
rect 126 32678 900 32684
rect 1548 32684 1554 32687
rect 1548 32678 1584 32684
rect 126 32644 138 32678
rect 1572 32644 1584 32678
rect 126 32638 900 32644
rect 894 32635 900 32638
rect 1548 32638 1584 32644
rect 1548 32635 1554 32638
rect 156 32598 162 32601
rect 126 32592 162 32598
rect 810 32598 816 32601
rect 810 32592 1584 32598
rect 126 32558 138 32592
rect 1572 32558 1584 32592
rect 126 32552 162 32558
rect 156 32549 162 32552
rect 810 32552 1584 32558
rect 810 32549 816 32552
rect 894 32512 900 32515
rect 126 32506 900 32512
rect 1548 32512 1554 32515
rect 1548 32506 1584 32512
rect 126 32472 138 32506
rect 1572 32472 1584 32506
rect 126 32466 900 32472
rect 894 32463 900 32466
rect 1548 32466 1584 32472
rect 1548 32463 1554 32466
rect 156 32426 162 32429
rect 126 32420 162 32426
rect 810 32426 816 32429
rect 810 32420 1584 32426
rect 126 32386 138 32420
rect 1572 32386 1584 32420
rect 126 32380 162 32386
rect 156 32377 162 32380
rect 810 32380 1584 32386
rect 810 32377 816 32380
rect 894 32340 900 32343
rect 126 32334 900 32340
rect 1548 32340 1554 32343
rect 1548 32334 1584 32340
rect 126 32300 138 32334
rect 1572 32300 1584 32334
rect 126 32294 900 32300
rect 894 32291 900 32294
rect 1548 32294 1584 32300
rect 1548 32291 1554 32294
rect 156 32254 162 32257
rect 126 32248 162 32254
rect 810 32254 816 32257
rect 810 32248 1584 32254
rect 126 32214 138 32248
rect 1572 32214 1584 32248
rect 126 32208 162 32214
rect 156 32205 162 32208
rect 810 32208 1584 32214
rect 810 32205 816 32208
rect 894 32168 900 32171
rect 126 32162 900 32168
rect 1548 32168 1554 32171
rect 1548 32162 1584 32168
rect 126 32128 138 32162
rect 1572 32128 1584 32162
rect 126 32122 900 32128
rect 894 32119 900 32122
rect 1548 32122 1584 32128
rect 1548 32119 1554 32122
rect 156 32082 162 32085
rect 126 32076 162 32082
rect 810 32082 816 32085
rect 810 32076 1584 32082
rect 126 32042 138 32076
rect 1572 32042 1584 32076
rect 126 32036 162 32042
rect 156 32033 162 32036
rect 810 32036 1584 32042
rect 810 32033 816 32036
rect 894 31996 900 31999
rect 126 31990 900 31996
rect 1548 31996 1554 31999
rect 1548 31990 1584 31996
rect 126 31956 138 31990
rect 1572 31956 1584 31990
rect 126 31950 900 31956
rect 894 31947 900 31950
rect 1548 31950 1584 31956
rect 1548 31947 1554 31950
rect 156 31910 162 31913
rect 126 31904 162 31910
rect 810 31910 816 31913
rect 810 31904 1584 31910
rect 126 31870 138 31904
rect 1572 31870 1584 31904
rect 126 31864 162 31870
rect 156 31861 162 31864
rect 810 31864 1584 31870
rect 810 31861 816 31864
rect 894 31824 900 31827
rect 126 31818 900 31824
rect 1548 31824 1554 31827
rect 1548 31818 1584 31824
rect 126 31784 138 31818
rect 1572 31784 1584 31818
rect 126 31778 900 31784
rect 894 31775 900 31778
rect 1548 31778 1584 31784
rect 1548 31775 1554 31778
rect 156 31738 162 31741
rect 126 31732 162 31738
rect 810 31738 816 31741
rect 810 31732 1584 31738
rect 126 31698 138 31732
rect 1572 31698 1584 31732
rect 126 31692 162 31698
rect 156 31689 162 31692
rect 810 31692 1584 31698
rect 810 31689 816 31692
rect 894 31652 900 31655
rect 126 31646 900 31652
rect 1548 31652 1554 31655
rect 1548 31646 1584 31652
rect 126 31612 138 31646
rect 1572 31612 1584 31646
rect 126 31606 900 31612
rect 894 31603 900 31606
rect 1548 31606 1584 31612
rect 1548 31603 1554 31606
rect 156 31566 162 31569
rect 126 31560 162 31566
rect 810 31566 816 31569
rect 810 31560 1584 31566
rect 126 31526 138 31560
rect 1572 31526 1584 31560
rect 126 31520 162 31526
rect 156 31517 162 31520
rect 810 31520 1584 31526
rect 810 31517 816 31520
rect 894 31480 900 31483
rect 126 31474 900 31480
rect 1548 31480 1554 31483
rect 1548 31474 1584 31480
rect 126 31440 138 31474
rect 1572 31440 1584 31474
rect 126 31434 900 31440
rect 894 31431 900 31434
rect 1548 31434 1584 31440
rect 1548 31431 1554 31434
rect 156 31394 162 31397
rect 126 31388 162 31394
rect 810 31394 816 31397
rect 810 31388 1584 31394
rect 126 31354 138 31388
rect 1572 31354 1584 31388
rect 126 31348 162 31354
rect 156 31345 162 31348
rect 810 31348 1584 31354
rect 810 31345 816 31348
rect 894 31308 900 31311
rect 126 31302 900 31308
rect 1548 31308 1554 31311
rect 1548 31302 1584 31308
rect 126 31268 138 31302
rect 1572 31268 1584 31302
rect 126 31262 900 31268
rect 894 31259 900 31262
rect 1548 31262 1584 31268
rect 1548 31259 1554 31262
rect 156 31222 162 31225
rect 126 31216 162 31222
rect 810 31222 816 31225
rect 810 31216 1584 31222
rect 126 31182 138 31216
rect 1572 31182 1584 31216
rect 126 31176 162 31182
rect 156 31173 162 31176
rect 810 31176 1584 31182
rect 810 31173 816 31176
rect 894 31136 900 31139
rect 126 31130 900 31136
rect 1548 31136 1554 31139
rect 1548 31130 1584 31136
rect 126 31096 138 31130
rect 1572 31096 1584 31130
rect 126 31090 900 31096
rect 894 31087 900 31090
rect 1548 31090 1584 31096
rect 1548 31087 1554 31090
rect 156 31050 162 31053
rect 126 31044 162 31050
rect 810 31050 816 31053
rect 810 31044 1584 31050
rect 126 31010 138 31044
rect 1572 31010 1584 31044
rect 126 31004 162 31010
rect 156 31001 162 31004
rect 810 31004 1584 31010
rect 810 31001 816 31004
rect 894 30964 900 30967
rect 126 30958 900 30964
rect 1548 30964 1554 30967
rect 1548 30958 1584 30964
rect 126 30924 138 30958
rect 1572 30924 1584 30958
rect 126 30918 900 30924
rect 894 30915 900 30918
rect 1548 30918 1584 30924
rect 1548 30915 1554 30918
rect 156 30878 162 30881
rect 126 30872 162 30878
rect 810 30878 816 30881
rect 810 30872 1584 30878
rect 126 30838 138 30872
rect 1572 30838 1584 30872
rect 126 30832 162 30838
rect 156 30829 162 30832
rect 810 30832 1584 30838
rect 810 30829 816 30832
rect 894 30792 900 30795
rect 126 30786 900 30792
rect 1548 30792 1554 30795
rect 1548 30786 1584 30792
rect 126 30752 138 30786
rect 1572 30752 1584 30786
rect 126 30746 900 30752
rect 894 30743 900 30746
rect 1548 30746 1584 30752
rect 1548 30743 1554 30746
rect 156 30706 162 30709
rect 126 30700 162 30706
rect 810 30706 816 30709
rect 810 30700 1584 30706
rect 126 30666 138 30700
rect 1572 30666 1584 30700
rect 126 30660 162 30666
rect 156 30657 162 30660
rect 810 30660 1584 30666
rect 810 30657 816 30660
rect 894 30620 900 30623
rect 126 30614 900 30620
rect 1548 30620 1554 30623
rect 1548 30614 1584 30620
rect 126 30580 138 30614
rect 1572 30580 1584 30614
rect 126 30574 900 30580
rect 894 30571 900 30574
rect 1548 30574 1584 30580
rect 1548 30571 1554 30574
rect 156 30534 162 30537
rect 126 30528 162 30534
rect 810 30534 816 30537
rect 810 30528 1584 30534
rect 126 30494 138 30528
rect 1572 30494 1584 30528
rect 126 30488 162 30494
rect 156 30485 162 30488
rect 810 30488 1584 30494
rect 810 30485 816 30488
rect 894 30448 900 30451
rect 126 30442 900 30448
rect 1548 30448 1554 30451
rect 1548 30442 1584 30448
rect 126 30408 138 30442
rect 1572 30408 1584 30442
rect 126 30402 900 30408
rect 894 30399 900 30402
rect 1548 30402 1584 30408
rect 1548 30399 1554 30402
rect 156 30362 162 30365
rect 126 30356 162 30362
rect 810 30362 816 30365
rect 810 30356 1584 30362
rect 126 30322 138 30356
rect 1572 30322 1584 30356
rect 126 30316 162 30322
rect 156 30313 162 30316
rect 810 30316 1584 30322
rect 810 30313 816 30316
rect 894 30276 900 30279
rect 126 30270 900 30276
rect 1548 30276 1554 30279
rect 1548 30270 1584 30276
rect 126 30236 138 30270
rect 1572 30236 1584 30270
rect 126 30230 900 30236
rect 894 30227 900 30230
rect 1548 30230 1584 30236
rect 1548 30227 1554 30230
rect 156 30190 162 30193
rect 126 30184 162 30190
rect 810 30190 816 30193
rect 810 30184 1584 30190
rect 126 30150 138 30184
rect 1572 30150 1584 30184
rect 126 30144 162 30150
rect 156 30141 162 30144
rect 810 30144 1584 30150
rect 810 30141 816 30144
rect 894 30104 900 30107
rect 126 30098 900 30104
rect 1548 30104 1554 30107
rect 1548 30098 1584 30104
rect 126 30064 138 30098
rect 1572 30064 1584 30098
rect 126 30058 900 30064
rect 894 30055 900 30058
rect 1548 30058 1584 30064
rect 1548 30055 1554 30058
rect 156 30018 162 30021
rect 126 30012 162 30018
rect 810 30018 816 30021
rect 810 30012 1584 30018
rect 126 29978 138 30012
rect 1572 29978 1584 30012
rect 126 29972 162 29978
rect 156 29969 162 29972
rect 810 29972 1584 29978
rect 810 29969 816 29972
rect 894 29932 900 29935
rect 126 29926 900 29932
rect 1548 29932 1554 29935
rect 1548 29926 1584 29932
rect 126 29892 138 29926
rect 1572 29892 1584 29926
rect 126 29886 900 29892
rect 894 29883 900 29886
rect 1548 29886 1584 29892
rect 1548 29883 1554 29886
rect 156 29846 162 29849
rect 126 29840 162 29846
rect 810 29846 816 29849
rect 810 29840 1584 29846
rect 126 29806 138 29840
rect 1572 29806 1584 29840
rect 126 29800 162 29806
rect 156 29797 162 29800
rect 810 29800 1584 29806
rect 810 29797 816 29800
rect 894 29760 900 29763
rect 126 29754 900 29760
rect 1548 29760 1554 29763
rect 1548 29754 1584 29760
rect 126 29720 138 29754
rect 1572 29720 1584 29754
rect 126 29714 900 29720
rect 894 29711 900 29714
rect 1548 29714 1584 29720
rect 1548 29711 1554 29714
rect 156 29674 162 29677
rect 126 29668 162 29674
rect 810 29674 816 29677
rect 810 29668 1584 29674
rect 126 29634 138 29668
rect 1572 29634 1584 29668
rect 126 29628 162 29634
rect 156 29625 162 29628
rect 810 29628 1584 29634
rect 810 29625 816 29628
rect 894 29588 900 29591
rect 126 29582 900 29588
rect 1548 29588 1554 29591
rect 1548 29582 1584 29588
rect 126 29548 138 29582
rect 1572 29548 1584 29582
rect 126 29542 900 29548
rect 894 29539 900 29542
rect 1548 29542 1584 29548
rect 1548 29539 1554 29542
rect 156 29502 162 29505
rect 126 29496 162 29502
rect 810 29502 816 29505
rect 810 29496 1584 29502
rect 126 29462 138 29496
rect 1572 29462 1584 29496
rect 126 29456 162 29462
rect 156 29453 162 29456
rect 810 29456 1584 29462
rect 810 29453 816 29456
rect 894 29416 900 29419
rect 126 29410 900 29416
rect 1548 29416 1554 29419
rect 1548 29410 1584 29416
rect 126 29376 138 29410
rect 1572 29376 1584 29410
rect 126 29370 900 29376
rect 894 29367 900 29370
rect 1548 29370 1584 29376
rect 1548 29367 1554 29370
rect 156 29330 162 29333
rect 126 29324 162 29330
rect 810 29330 816 29333
rect 810 29324 1584 29330
rect 126 29290 138 29324
rect 1572 29290 1584 29324
rect 126 29284 162 29290
rect 156 29281 162 29284
rect 810 29284 1584 29290
rect 810 29281 816 29284
rect 894 29244 900 29247
rect 126 29238 900 29244
rect 1548 29244 1554 29247
rect 1548 29238 1584 29244
rect 126 29204 138 29238
rect 1572 29204 1584 29238
rect 126 29198 900 29204
rect 894 29195 900 29198
rect 1548 29198 1584 29204
rect 1548 29195 1554 29198
rect 156 29158 162 29161
rect 126 29152 162 29158
rect 810 29158 816 29161
rect 810 29152 1584 29158
rect 126 29118 138 29152
rect 1572 29118 1584 29152
rect 126 29112 162 29118
rect 156 29109 162 29112
rect 810 29112 1584 29118
rect 810 29109 816 29112
rect 894 29072 900 29075
rect 126 29066 900 29072
rect 1548 29072 1554 29075
rect 1548 29066 1584 29072
rect 126 29032 138 29066
rect 1572 29032 1584 29066
rect 126 29026 900 29032
rect 894 29023 900 29026
rect 1548 29026 1584 29032
rect 1548 29023 1554 29026
rect 156 28986 162 28989
rect 126 28980 162 28986
rect 810 28986 816 28989
rect 810 28980 1584 28986
rect 126 28946 138 28980
rect 1572 28946 1584 28980
rect 126 28940 162 28946
rect 156 28937 162 28940
rect 810 28940 1584 28946
rect 810 28937 816 28940
rect 894 28900 900 28903
rect 126 28894 900 28900
rect 1548 28900 1554 28903
rect 1548 28894 1584 28900
rect 126 28860 138 28894
rect 1572 28860 1584 28894
rect 126 28854 900 28860
rect 894 28851 900 28854
rect 1548 28854 1584 28860
rect 1548 28851 1554 28854
rect 156 28814 162 28817
rect 126 28808 162 28814
rect 810 28814 816 28817
rect 810 28808 1584 28814
rect 126 28774 138 28808
rect 1572 28774 1584 28808
rect 126 28768 162 28774
rect 156 28765 162 28768
rect 810 28768 1584 28774
rect 810 28765 816 28768
rect 894 28728 900 28731
rect 126 28722 900 28728
rect 1548 28728 1554 28731
rect 1548 28722 1584 28728
rect 126 28688 138 28722
rect 1572 28688 1584 28722
rect 126 28682 900 28688
rect 894 28679 900 28682
rect 1548 28682 1584 28688
rect 1548 28679 1554 28682
rect 156 28642 162 28645
rect 126 28636 162 28642
rect 810 28642 816 28645
rect 810 28636 1584 28642
rect 126 28602 138 28636
rect 1572 28602 1584 28636
rect 126 28596 162 28602
rect 156 28593 162 28596
rect 810 28596 1584 28602
rect 810 28593 816 28596
rect 894 28556 900 28559
rect 126 28550 900 28556
rect 1548 28556 1554 28559
rect 1548 28550 1584 28556
rect 126 28516 138 28550
rect 1572 28516 1584 28550
rect 126 28510 900 28516
rect 894 28507 900 28510
rect 1548 28510 1584 28516
rect 1548 28507 1554 28510
rect 156 28470 162 28473
rect 126 28464 162 28470
rect 810 28470 816 28473
rect 810 28464 1584 28470
rect 126 28430 138 28464
rect 1572 28430 1584 28464
rect 126 28424 162 28430
rect 156 28421 162 28424
rect 810 28424 1584 28430
rect 810 28421 816 28424
rect 894 28384 900 28387
rect 126 28378 900 28384
rect 1548 28384 1554 28387
rect 1548 28378 1584 28384
rect 126 28344 138 28378
rect 1572 28344 1584 28378
rect 126 28338 900 28344
rect 894 28335 900 28338
rect 1548 28338 1584 28344
rect 1548 28335 1554 28338
rect 156 28298 162 28301
rect 126 28292 162 28298
rect 810 28298 816 28301
rect 810 28292 1584 28298
rect 126 28258 138 28292
rect 1572 28258 1584 28292
rect 126 28252 162 28258
rect 156 28249 162 28252
rect 810 28252 1584 28258
rect 810 28249 816 28252
rect 894 28212 900 28215
rect 126 28206 900 28212
rect 1548 28212 1554 28215
rect 1548 28206 1584 28212
rect 126 28172 138 28206
rect 1572 28172 1584 28206
rect 126 28166 900 28172
rect 894 28163 900 28166
rect 1548 28166 1584 28172
rect 1548 28163 1554 28166
rect 156 28126 162 28129
rect 126 28120 162 28126
rect 810 28126 816 28129
rect 810 28120 1584 28126
rect 126 28086 138 28120
rect 1572 28086 1584 28120
rect 126 28080 162 28086
rect 156 28077 162 28080
rect 810 28080 1584 28086
rect 810 28077 816 28080
rect 894 28040 900 28043
rect 126 28034 900 28040
rect 1548 28040 1554 28043
rect 1548 28034 1584 28040
rect 126 28000 138 28034
rect 1572 28000 1584 28034
rect 126 27994 900 28000
rect 894 27991 900 27994
rect 1548 27994 1584 28000
rect 1548 27991 1554 27994
rect 156 27954 162 27957
rect 126 27948 162 27954
rect 810 27954 816 27957
rect 810 27948 1584 27954
rect 126 27914 138 27948
rect 1572 27914 1584 27948
rect 126 27908 162 27914
rect 156 27905 162 27908
rect 810 27908 1584 27914
rect 810 27905 816 27908
rect 894 27868 900 27871
rect 126 27862 900 27868
rect 1548 27868 1554 27871
rect 1548 27862 1584 27868
rect 126 27828 138 27862
rect 1572 27828 1584 27862
rect 126 27822 900 27828
rect 894 27819 900 27822
rect 1548 27822 1584 27828
rect 1548 27819 1554 27822
rect 156 27782 162 27785
rect 126 27776 162 27782
rect 810 27782 816 27785
rect 810 27776 1584 27782
rect 126 27742 138 27776
rect 1572 27742 1584 27776
rect 126 27736 162 27742
rect 156 27733 162 27736
rect 810 27736 1584 27742
rect 810 27733 816 27736
rect 894 27696 900 27699
rect 126 27690 900 27696
rect 1548 27696 1554 27699
rect 1548 27690 1584 27696
rect 126 27656 138 27690
rect 1572 27656 1584 27690
rect 126 27650 900 27656
rect 894 27647 900 27650
rect 1548 27650 1584 27656
rect 1548 27647 1554 27650
rect 156 27610 162 27613
rect 126 27604 162 27610
rect 810 27610 816 27613
rect 810 27604 1584 27610
rect 126 27570 138 27604
rect 1572 27570 1584 27604
rect 126 27564 162 27570
rect 156 27561 162 27564
rect 810 27564 1584 27570
rect 810 27561 816 27564
rect 894 27524 900 27527
rect 126 27518 900 27524
rect 1548 27524 1554 27527
rect 1548 27518 1584 27524
rect 126 27484 138 27518
rect 1572 27484 1584 27518
rect 126 27478 900 27484
rect 894 27475 900 27478
rect 1548 27478 1584 27484
rect 1548 27475 1554 27478
rect 156 27438 162 27441
rect 126 27432 162 27438
rect 810 27438 816 27441
rect 810 27432 1584 27438
rect 126 27398 138 27432
rect 1572 27398 1584 27432
rect 126 27392 162 27398
rect 156 27389 162 27392
rect 810 27392 1584 27398
rect 810 27389 816 27392
rect 894 27352 900 27355
rect 126 27346 900 27352
rect 1548 27352 1554 27355
rect 1548 27346 1584 27352
rect 126 27312 138 27346
rect 1572 27312 1584 27346
rect 126 27306 900 27312
rect 894 27303 900 27306
rect 1548 27306 1584 27312
rect 1548 27303 1554 27306
rect 156 27266 162 27269
rect 126 27260 162 27266
rect 810 27266 816 27269
rect 810 27260 1584 27266
rect 126 27226 138 27260
rect 1572 27226 1584 27260
rect 126 27220 162 27226
rect 156 27217 162 27220
rect 810 27220 1584 27226
rect 810 27217 816 27220
rect 894 27180 900 27183
rect 126 27174 900 27180
rect 1548 27180 1554 27183
rect 1548 27174 1584 27180
rect 126 27140 138 27174
rect 1572 27140 1584 27174
rect 126 27134 900 27140
rect 894 27131 900 27134
rect 1548 27134 1584 27140
rect 1548 27131 1554 27134
rect 156 27094 162 27097
rect 126 27088 162 27094
rect 810 27094 816 27097
rect 810 27088 1584 27094
rect 126 27054 138 27088
rect 1572 27054 1584 27088
rect 126 27048 162 27054
rect 156 27045 162 27048
rect 810 27048 1584 27054
rect 810 27045 816 27048
rect 894 27008 900 27011
rect 126 27002 900 27008
rect 1548 27008 1554 27011
rect 1548 27002 1584 27008
rect 126 26968 138 27002
rect 1572 26968 1584 27002
rect 126 26962 900 26968
rect 894 26959 900 26962
rect 1548 26962 1584 26968
rect 1548 26959 1554 26962
rect 156 26922 162 26925
rect 126 26916 162 26922
rect 810 26922 816 26925
rect 810 26916 1584 26922
rect 126 26882 138 26916
rect 1572 26882 1584 26916
rect 126 26876 162 26882
rect 156 26873 162 26876
rect 810 26876 1584 26882
rect 810 26873 816 26876
rect 894 26836 900 26839
rect 126 26830 900 26836
rect 1548 26836 1554 26839
rect 1548 26830 1584 26836
rect 126 26796 138 26830
rect 1572 26796 1584 26830
rect 126 26790 900 26796
rect 894 26787 900 26790
rect 1548 26790 1584 26796
rect 1548 26787 1554 26790
rect 156 26750 162 26753
rect 126 26744 162 26750
rect 810 26750 816 26753
rect 810 26744 1584 26750
rect 126 26710 138 26744
rect 1572 26710 1584 26744
rect 126 26704 162 26710
rect 156 26701 162 26704
rect 810 26704 1584 26710
rect 810 26701 816 26704
rect 894 26664 900 26667
rect 126 26658 900 26664
rect 1548 26664 1554 26667
rect 1548 26658 1584 26664
rect 126 26624 138 26658
rect 1572 26624 1584 26658
rect 126 26618 900 26624
rect 894 26615 900 26618
rect 1548 26618 1584 26624
rect 1548 26615 1554 26618
rect 156 26578 162 26581
rect 126 26572 162 26578
rect 810 26578 816 26581
rect 810 26572 1584 26578
rect 126 26538 138 26572
rect 1572 26538 1584 26572
rect 126 26532 162 26538
rect 156 26529 162 26532
rect 810 26532 1584 26538
rect 810 26529 816 26532
rect 894 26492 900 26495
rect 126 26486 900 26492
rect 1548 26492 1554 26495
rect 1548 26486 1584 26492
rect 126 26452 138 26486
rect 1572 26452 1584 26486
rect 126 26446 900 26452
rect 894 26443 900 26446
rect 1548 26446 1584 26452
rect 1548 26443 1554 26446
rect 156 26406 162 26409
rect 126 26400 162 26406
rect 810 26406 816 26409
rect 810 26400 1584 26406
rect 126 26366 138 26400
rect 1572 26366 1584 26400
rect 126 26360 162 26366
rect 156 26357 162 26360
rect 810 26360 1584 26366
rect 810 26357 816 26360
rect 894 26320 900 26323
rect 126 26314 900 26320
rect 1548 26320 1554 26323
rect 1548 26314 1584 26320
rect 126 26280 138 26314
rect 1572 26280 1584 26314
rect 126 26274 900 26280
rect 894 26271 900 26274
rect 1548 26274 1584 26280
rect 1548 26271 1554 26274
rect 156 26234 162 26237
rect 126 26228 162 26234
rect 810 26234 816 26237
rect 810 26228 1584 26234
rect 126 26194 138 26228
rect 1572 26194 1584 26228
rect 126 26188 162 26194
rect 156 26185 162 26188
rect 810 26188 1584 26194
rect 810 26185 816 26188
rect 894 26148 900 26151
rect 126 26142 900 26148
rect 1548 26148 1554 26151
rect 1548 26142 1584 26148
rect 126 26108 138 26142
rect 1572 26108 1584 26142
rect 126 26102 900 26108
rect 894 26099 900 26102
rect 1548 26102 1584 26108
rect 1548 26099 1554 26102
rect 156 26062 162 26065
rect 126 26056 162 26062
rect 810 26062 816 26065
rect 810 26056 1584 26062
rect 126 26022 138 26056
rect 1572 26022 1584 26056
rect 126 26016 162 26022
rect 156 26013 162 26016
rect 810 26016 1584 26022
rect 810 26013 816 26016
rect 894 25976 900 25979
rect 126 25970 900 25976
rect 1548 25976 1554 25979
rect 1548 25970 1584 25976
rect 126 25936 138 25970
rect 1572 25936 1584 25970
rect 126 25930 900 25936
rect 894 25927 900 25930
rect 1548 25930 1584 25936
rect 1548 25927 1554 25930
rect 156 25890 162 25893
rect 126 25884 162 25890
rect 810 25890 816 25893
rect 810 25884 1584 25890
rect 126 25850 138 25884
rect 1572 25850 1584 25884
rect 126 25844 162 25850
rect 156 25841 162 25844
rect 810 25844 1584 25850
rect 810 25841 816 25844
rect 894 25804 900 25807
rect 126 25798 900 25804
rect 1548 25804 1554 25807
rect 1548 25798 1584 25804
rect 126 25764 138 25798
rect 1572 25764 1584 25798
rect 126 25758 900 25764
rect 894 25755 900 25758
rect 1548 25758 1584 25764
rect 1548 25755 1554 25758
rect 156 25718 162 25721
rect 126 25712 162 25718
rect 810 25718 816 25721
rect 810 25712 1584 25718
rect 126 25678 138 25712
rect 1572 25678 1584 25712
rect 126 25672 162 25678
rect 156 25669 162 25672
rect 810 25672 1584 25678
rect 810 25669 816 25672
rect 894 25632 900 25635
rect 126 25626 900 25632
rect 1548 25632 1554 25635
rect 1548 25626 1584 25632
rect 126 25592 138 25626
rect 1572 25592 1584 25626
rect 126 25586 900 25592
rect 894 25583 900 25586
rect 1548 25586 1584 25592
rect 1548 25583 1554 25586
rect 156 25546 162 25549
rect 126 25540 162 25546
rect 810 25546 816 25549
rect 810 25540 1584 25546
rect 126 25506 138 25540
rect 1572 25506 1584 25540
rect 126 25500 162 25506
rect 156 25497 162 25500
rect 810 25500 1584 25506
rect 810 25497 816 25500
rect 894 25460 900 25463
rect 126 25454 900 25460
rect 1548 25460 1554 25463
rect 1548 25454 1584 25460
rect 126 25420 138 25454
rect 1572 25420 1584 25454
rect 126 25414 900 25420
rect 894 25411 900 25414
rect 1548 25414 1584 25420
rect 1548 25411 1554 25414
rect 156 25374 162 25377
rect 126 25368 162 25374
rect 810 25374 816 25377
rect 810 25368 1584 25374
rect 126 25334 138 25368
rect 1572 25334 1584 25368
rect 126 25328 162 25334
rect 156 25325 162 25328
rect 810 25328 1584 25334
rect 810 25325 816 25328
rect 894 25288 900 25291
rect 126 25282 900 25288
rect 1548 25288 1554 25291
rect 1548 25282 1584 25288
rect 126 25248 138 25282
rect 1572 25248 1584 25282
rect 126 25242 900 25248
rect 894 25239 900 25242
rect 1548 25242 1584 25248
rect 1548 25239 1554 25242
rect 156 25202 162 25205
rect 126 25196 162 25202
rect 810 25202 816 25205
rect 810 25196 1584 25202
rect 126 25162 138 25196
rect 1572 25162 1584 25196
rect 126 25156 162 25162
rect 156 25153 162 25156
rect 810 25156 1584 25162
rect 810 25153 816 25156
rect 894 25116 900 25119
rect 126 25110 900 25116
rect 1548 25116 1554 25119
rect 1548 25110 1584 25116
rect 126 25076 138 25110
rect 1572 25076 1584 25110
rect 126 25070 900 25076
rect 894 25067 900 25070
rect 1548 25070 1584 25076
rect 1548 25067 1554 25070
rect 156 25030 162 25033
rect 126 25024 162 25030
rect 810 25030 816 25033
rect 810 25024 1584 25030
rect 126 24990 138 25024
rect 1572 24990 1584 25024
rect 126 24984 162 24990
rect 156 24981 162 24984
rect 810 24984 1584 24990
rect 810 24981 816 24984
rect 894 24944 900 24947
rect 126 24938 900 24944
rect 1548 24944 1554 24947
rect 1548 24938 1584 24944
rect 126 24904 138 24938
rect 1572 24904 1584 24938
rect 126 24898 900 24904
rect 894 24895 900 24898
rect 1548 24898 1584 24904
rect 1548 24895 1554 24898
rect 156 24858 162 24861
rect 126 24852 162 24858
rect 810 24858 816 24861
rect 810 24852 1584 24858
rect 126 24818 138 24852
rect 1572 24818 1584 24852
rect 126 24812 162 24818
rect 156 24809 162 24812
rect 810 24812 1584 24818
rect 810 24809 816 24812
rect 894 24772 900 24775
rect 126 24766 900 24772
rect 1548 24772 1554 24775
rect 1548 24766 1584 24772
rect 126 24732 138 24766
rect 1572 24732 1584 24766
rect 126 24726 900 24732
rect 894 24723 900 24726
rect 1548 24726 1584 24732
rect 1548 24723 1554 24726
rect 156 24686 162 24689
rect 126 24680 162 24686
rect 810 24686 816 24689
rect 810 24680 1584 24686
rect 126 24646 138 24680
rect 1572 24646 1584 24680
rect 126 24640 162 24646
rect 156 24637 162 24640
rect 810 24640 1584 24646
rect 810 24637 816 24640
rect 894 24600 900 24603
rect 126 24594 900 24600
rect 1548 24600 1554 24603
rect 1548 24594 1584 24600
rect 126 24560 138 24594
rect 1572 24560 1584 24594
rect 126 24554 900 24560
rect 894 24551 900 24554
rect 1548 24554 1584 24560
rect 1548 24551 1554 24554
rect 156 24514 162 24517
rect 126 24508 162 24514
rect 810 24514 816 24517
rect 810 24508 1584 24514
rect 126 24474 138 24508
rect 1572 24474 1584 24508
rect 126 24468 162 24474
rect 156 24465 162 24468
rect 810 24468 1584 24474
rect 810 24465 816 24468
rect 894 24428 900 24431
rect 126 24422 900 24428
rect 1548 24428 1554 24431
rect 1548 24422 1584 24428
rect 126 24388 138 24422
rect 1572 24388 1584 24422
rect 126 24382 900 24388
rect 894 24379 900 24382
rect 1548 24382 1584 24388
rect 1548 24379 1554 24382
rect 156 24342 162 24345
rect 126 24336 162 24342
rect 810 24342 816 24345
rect 810 24336 1584 24342
rect 126 24302 138 24336
rect 1572 24302 1584 24336
rect 126 24296 162 24302
rect 156 24293 162 24296
rect 810 24296 1584 24302
rect 810 24293 816 24296
rect 894 24256 900 24259
rect 126 24250 900 24256
rect 1548 24256 1554 24259
rect 1548 24250 1584 24256
rect 126 24216 138 24250
rect 1572 24216 1584 24250
rect 126 24210 900 24216
rect 894 24207 900 24210
rect 1548 24210 1584 24216
rect 1548 24207 1554 24210
rect 156 24170 162 24173
rect 126 24164 162 24170
rect 810 24170 816 24173
rect 810 24164 1584 24170
rect 126 24130 138 24164
rect 1572 24130 1584 24164
rect 126 24124 162 24130
rect 156 24121 162 24124
rect 810 24124 1584 24130
rect 810 24121 816 24124
rect 894 24084 900 24087
rect 126 24078 900 24084
rect 1548 24084 1554 24087
rect 1548 24078 1584 24084
rect 126 24044 138 24078
rect 1572 24044 1584 24078
rect 126 24038 900 24044
rect 894 24035 900 24038
rect 1548 24038 1584 24044
rect 1548 24035 1554 24038
rect 156 23998 162 24001
rect 126 23992 162 23998
rect 810 23998 816 24001
rect 810 23992 1584 23998
rect 126 23958 138 23992
rect 1572 23958 1584 23992
rect 126 23952 162 23958
rect 156 23949 162 23952
rect 810 23952 1584 23958
rect 810 23949 816 23952
rect 894 23912 900 23915
rect 126 23906 900 23912
rect 1548 23912 1554 23915
rect 1548 23906 1584 23912
rect 126 23872 138 23906
rect 1572 23872 1584 23906
rect 126 23866 900 23872
rect 894 23863 900 23866
rect 1548 23866 1584 23872
rect 1548 23863 1554 23866
rect 156 23826 162 23829
rect 126 23820 162 23826
rect 810 23826 816 23829
rect 810 23820 1584 23826
rect 126 23786 138 23820
rect 1572 23786 1584 23820
rect 126 23780 162 23786
rect 156 23777 162 23780
rect 810 23780 1584 23786
rect 810 23777 816 23780
rect 894 23740 900 23743
rect 126 23734 900 23740
rect 1548 23740 1554 23743
rect 1548 23734 1584 23740
rect 126 23700 138 23734
rect 1572 23700 1584 23734
rect 126 23694 900 23700
rect 894 23691 900 23694
rect 1548 23694 1584 23700
rect 1548 23691 1554 23694
rect 156 23654 162 23657
rect 126 23648 162 23654
rect 810 23654 816 23657
rect 810 23648 1584 23654
rect 126 23614 138 23648
rect 1572 23614 1584 23648
rect 126 23608 162 23614
rect 156 23605 162 23608
rect 810 23608 1584 23614
rect 810 23605 816 23608
rect 894 23568 900 23571
rect 126 23562 900 23568
rect 1548 23568 1554 23571
rect 1548 23562 1584 23568
rect 126 23528 138 23562
rect 1572 23528 1584 23562
rect 126 23522 900 23528
rect 894 23519 900 23522
rect 1548 23522 1584 23528
rect 1548 23519 1554 23522
rect 156 23482 162 23485
rect 126 23476 162 23482
rect 810 23482 816 23485
rect 810 23476 1584 23482
rect 126 23442 138 23476
rect 1572 23442 1584 23476
rect 126 23436 162 23442
rect 156 23433 162 23436
rect 810 23436 1584 23442
rect 810 23433 816 23436
rect 894 23396 900 23399
rect 126 23390 900 23396
rect 1548 23396 1554 23399
rect 1548 23390 1584 23396
rect 126 23356 138 23390
rect 1572 23356 1584 23390
rect 126 23350 900 23356
rect 894 23347 900 23350
rect 1548 23350 1584 23356
rect 1548 23347 1554 23350
rect 156 23310 162 23313
rect 126 23304 162 23310
rect 810 23310 816 23313
rect 810 23304 1584 23310
rect 126 23270 138 23304
rect 1572 23270 1584 23304
rect 126 23264 162 23270
rect 156 23261 162 23264
rect 810 23264 1584 23270
rect 810 23261 816 23264
rect 894 23224 900 23227
rect 126 23218 900 23224
rect 1548 23224 1554 23227
rect 1548 23218 1584 23224
rect 126 23184 138 23218
rect 1572 23184 1584 23218
rect 126 23178 900 23184
rect 894 23175 900 23178
rect 1548 23178 1584 23184
rect 1548 23175 1554 23178
rect 156 23138 162 23141
rect 126 23132 162 23138
rect 810 23138 816 23141
rect 810 23132 1584 23138
rect 126 23098 138 23132
rect 1572 23098 1584 23132
rect 126 23092 162 23098
rect 156 23089 162 23092
rect 810 23092 1584 23098
rect 810 23089 816 23092
rect 894 23052 900 23055
rect 126 23046 900 23052
rect 1548 23052 1554 23055
rect 1548 23046 1584 23052
rect 126 23012 138 23046
rect 1572 23012 1584 23046
rect 126 23006 900 23012
rect 894 23003 900 23006
rect 1548 23006 1584 23012
rect 1548 23003 1554 23006
rect 156 22966 162 22969
rect 126 22960 162 22966
rect 810 22966 816 22969
rect 810 22960 1584 22966
rect 126 22926 138 22960
rect 1572 22926 1584 22960
rect 126 22920 162 22926
rect 156 22917 162 22920
rect 810 22920 1584 22926
rect 810 22917 816 22920
rect 894 22880 900 22883
rect 126 22874 900 22880
rect 1548 22880 1554 22883
rect 1548 22874 1584 22880
rect 126 22840 138 22874
rect 1572 22840 1584 22874
rect 126 22834 900 22840
rect 894 22831 900 22834
rect 1548 22834 1584 22840
rect 1548 22831 1554 22834
rect 156 22794 162 22797
rect 126 22788 162 22794
rect 810 22794 816 22797
rect 810 22788 1584 22794
rect 126 22754 138 22788
rect 1572 22754 1584 22788
rect 126 22748 162 22754
rect 156 22745 162 22748
rect 810 22748 1584 22754
rect 810 22745 816 22748
rect 894 22708 900 22711
rect 126 22702 900 22708
rect 1548 22708 1554 22711
rect 1548 22702 1584 22708
rect 126 22668 138 22702
rect 1572 22668 1584 22702
rect 126 22662 900 22668
rect 894 22659 900 22662
rect 1548 22662 1584 22668
rect 1548 22659 1554 22662
rect 156 22622 162 22625
rect 126 22616 162 22622
rect 810 22622 816 22625
rect 810 22616 1584 22622
rect 126 22582 138 22616
rect 1572 22582 1584 22616
rect 126 22576 162 22582
rect 156 22573 162 22576
rect 810 22576 1584 22582
rect 810 22573 816 22576
rect 894 22536 900 22539
rect 126 22530 900 22536
rect 1548 22536 1554 22539
rect 1548 22530 1584 22536
rect 126 22496 138 22530
rect 1572 22496 1584 22530
rect 126 22490 900 22496
rect 894 22487 900 22490
rect 1548 22490 1584 22496
rect 1548 22487 1554 22490
rect 156 22450 162 22453
rect 126 22444 162 22450
rect 810 22450 816 22453
rect 810 22444 1584 22450
rect 126 22410 138 22444
rect 1572 22410 1584 22444
rect 126 22404 162 22410
rect 156 22401 162 22404
rect 810 22404 1584 22410
rect 810 22401 816 22404
rect 894 22364 900 22367
rect 126 22358 900 22364
rect 1548 22364 1554 22367
rect 1548 22358 1584 22364
rect 126 22324 138 22358
rect 1572 22324 1584 22358
rect 126 22318 900 22324
rect 894 22315 900 22318
rect 1548 22318 1584 22324
rect 1548 22315 1554 22318
rect 156 22278 162 22281
rect 126 22272 162 22278
rect 810 22278 816 22281
rect 810 22272 1584 22278
rect 126 22238 138 22272
rect 1572 22238 1584 22272
rect 126 22232 162 22238
rect 156 22229 162 22232
rect 810 22232 1584 22238
rect 810 22229 816 22232
rect 894 22192 900 22195
rect 126 22186 900 22192
rect 1548 22192 1554 22195
rect 1548 22186 1584 22192
rect 126 22152 138 22186
rect 1572 22152 1584 22186
rect 126 22146 900 22152
rect 894 22143 900 22146
rect 1548 22146 1584 22152
rect 1548 22143 1554 22146
rect 156 22106 162 22109
rect 126 22100 162 22106
rect 810 22106 816 22109
rect 810 22100 1584 22106
rect 126 22066 138 22100
rect 1572 22066 1584 22100
rect 126 22060 162 22066
rect 156 22057 162 22060
rect 810 22060 1584 22066
rect 810 22057 816 22060
rect 894 22020 900 22023
rect 126 22014 900 22020
rect 1548 22020 1554 22023
rect 1548 22014 1584 22020
rect 126 21980 138 22014
rect 1572 21980 1584 22014
rect 126 21974 900 21980
rect 894 21971 900 21974
rect 1548 21974 1584 21980
rect 1548 21971 1554 21974
rect 156 21934 162 21937
rect 126 21928 162 21934
rect 810 21934 816 21937
rect 810 21928 1584 21934
rect 126 21894 138 21928
rect 1572 21894 1584 21928
rect 126 21888 162 21894
rect 156 21885 162 21888
rect 810 21888 1584 21894
rect 810 21885 816 21888
rect 894 21848 900 21851
rect 126 21842 900 21848
rect 1548 21848 1554 21851
rect 1548 21842 1584 21848
rect 126 21808 138 21842
rect 1572 21808 1584 21842
rect 126 21802 900 21808
rect 894 21799 900 21802
rect 1548 21802 1584 21808
rect 1548 21799 1554 21802
rect 156 21762 162 21765
rect 126 21756 162 21762
rect 810 21762 816 21765
rect 810 21756 1584 21762
rect 126 21722 138 21756
rect 1572 21722 1584 21756
rect 126 21716 162 21722
rect 156 21713 162 21716
rect 810 21716 1584 21722
rect 810 21713 816 21716
rect 894 21676 900 21679
rect 126 21670 900 21676
rect 1548 21676 1554 21679
rect 1548 21670 1584 21676
rect 126 21636 138 21670
rect 1572 21636 1584 21670
rect 126 21630 900 21636
rect 894 21627 900 21630
rect 1548 21630 1584 21636
rect 1548 21627 1554 21630
rect 156 21590 162 21593
rect 126 21584 162 21590
rect 810 21590 816 21593
rect 810 21584 1584 21590
rect 126 21550 138 21584
rect 1572 21550 1584 21584
rect 126 21544 162 21550
rect 156 21541 162 21544
rect 810 21544 1584 21550
rect 810 21541 816 21544
rect 894 21504 900 21507
rect 126 21498 900 21504
rect 1548 21504 1554 21507
rect 1548 21498 1584 21504
rect 126 21464 138 21498
rect 1572 21464 1584 21498
rect 126 21458 900 21464
rect 894 21455 900 21458
rect 1548 21458 1584 21464
rect 1548 21455 1554 21458
rect 156 21418 162 21421
rect 126 21412 162 21418
rect 810 21418 816 21421
rect 810 21412 1584 21418
rect 126 21378 138 21412
rect 1572 21378 1584 21412
rect 126 21372 162 21378
rect 156 21369 162 21372
rect 810 21372 1584 21378
rect 810 21369 816 21372
rect 894 21332 900 21335
rect 126 21326 900 21332
rect 1548 21332 1554 21335
rect 1548 21326 1584 21332
rect 126 21292 138 21326
rect 1572 21292 1584 21326
rect 126 21286 900 21292
rect 894 21283 900 21286
rect 1548 21286 1584 21292
rect 1548 21283 1554 21286
rect 156 21246 162 21249
rect 126 21240 162 21246
rect 810 21246 816 21249
rect 810 21240 1584 21246
rect 126 21206 138 21240
rect 1572 21206 1584 21240
rect 126 21200 162 21206
rect 156 21197 162 21200
rect 810 21200 1584 21206
rect 810 21197 816 21200
rect 894 21160 900 21163
rect 126 21154 900 21160
rect 1548 21160 1554 21163
rect 1548 21154 1584 21160
rect 126 21120 138 21154
rect 1572 21120 1584 21154
rect 126 21114 900 21120
rect 894 21111 900 21114
rect 1548 21114 1584 21120
rect 1548 21111 1554 21114
rect 156 21074 162 21077
rect 126 21068 162 21074
rect 810 21074 816 21077
rect 810 21068 1584 21074
rect 126 21034 138 21068
rect 1572 21034 1584 21068
rect 126 21028 162 21034
rect 156 21025 162 21028
rect 810 21028 1584 21034
rect 810 21025 816 21028
rect 894 20988 900 20991
rect 126 20982 900 20988
rect 1548 20988 1554 20991
rect 1548 20982 1584 20988
rect 126 20948 138 20982
rect 1572 20948 1584 20982
rect 126 20942 900 20948
rect 894 20939 900 20942
rect 1548 20942 1584 20948
rect 1548 20939 1554 20942
rect 156 20902 162 20905
rect 126 20896 162 20902
rect 810 20902 816 20905
rect 810 20896 1584 20902
rect 126 20862 138 20896
rect 1572 20862 1584 20896
rect 126 20856 162 20862
rect 156 20853 162 20856
rect 810 20856 1584 20862
rect 810 20853 816 20856
rect 894 20816 900 20819
rect 126 20810 900 20816
rect 1548 20816 1554 20819
rect 1548 20810 1584 20816
rect 126 20776 138 20810
rect 1572 20776 1584 20810
rect 126 20770 900 20776
rect 894 20767 900 20770
rect 1548 20770 1584 20776
rect 1548 20767 1554 20770
rect 156 20730 162 20733
rect 126 20724 162 20730
rect 810 20730 816 20733
rect 810 20724 1584 20730
rect 126 20690 138 20724
rect 1572 20690 1584 20724
rect 126 20684 162 20690
rect 156 20681 162 20684
rect 810 20684 1584 20690
rect 810 20681 816 20684
rect 894 20644 900 20647
rect 126 20638 900 20644
rect 1548 20644 1554 20647
rect 1548 20638 1584 20644
rect 126 20604 138 20638
rect 1572 20604 1584 20638
rect 126 20598 900 20604
rect 894 20595 900 20598
rect 1548 20598 1584 20604
rect 1548 20595 1554 20598
rect 156 20558 162 20561
rect 126 20552 162 20558
rect 810 20558 816 20561
rect 810 20552 1584 20558
rect 126 20518 138 20552
rect 1572 20518 1584 20552
rect 126 20512 162 20518
rect 156 20509 162 20512
rect 810 20512 1584 20518
rect 810 20509 816 20512
rect 894 20472 900 20475
rect 126 20466 900 20472
rect 1548 20472 1554 20475
rect 1548 20466 1584 20472
rect 126 20432 138 20466
rect 1572 20432 1584 20466
rect 126 20426 900 20432
rect 894 20423 900 20426
rect 1548 20426 1584 20432
rect 1548 20423 1554 20426
rect 156 20386 162 20389
rect 126 20380 162 20386
rect 810 20386 816 20389
rect 810 20380 1584 20386
rect 126 20346 138 20380
rect 1572 20346 1584 20380
rect 126 20340 162 20346
rect 156 20337 162 20340
rect 810 20340 1584 20346
rect 810 20337 816 20340
rect 894 20300 900 20303
rect 126 20294 900 20300
rect 1548 20300 1554 20303
rect 1548 20294 1584 20300
rect 126 20260 138 20294
rect 1572 20260 1584 20294
rect 126 20254 900 20260
rect 894 20251 900 20254
rect 1548 20254 1584 20260
rect 1548 20251 1554 20254
rect 156 20214 162 20217
rect 126 20208 162 20214
rect 810 20214 816 20217
rect 810 20208 1584 20214
rect 126 20174 138 20208
rect 1572 20174 1584 20208
rect 126 20168 162 20174
rect 156 20165 162 20168
rect 810 20168 1584 20174
rect 810 20165 816 20168
rect 894 20128 900 20131
rect 126 20122 900 20128
rect 1548 20128 1554 20131
rect 1548 20122 1584 20128
rect 126 20088 138 20122
rect 1572 20088 1584 20122
rect 126 20082 900 20088
rect 894 20079 900 20082
rect 1548 20082 1584 20088
rect 1548 20079 1554 20082
rect 156 20042 162 20045
rect 126 20036 162 20042
rect 810 20042 816 20045
rect 810 20036 1584 20042
rect 126 20002 138 20036
rect 1572 20002 1584 20036
rect 126 19996 162 20002
rect 156 19993 162 19996
rect 810 19996 1584 20002
rect 810 19993 816 19996
rect 894 19956 900 19959
rect 126 19950 900 19956
rect 1548 19956 1554 19959
rect 1548 19950 1584 19956
rect 126 19916 138 19950
rect 1572 19916 1584 19950
rect 126 19910 900 19916
rect 894 19907 900 19910
rect 1548 19910 1584 19916
rect 1548 19907 1554 19910
rect 156 19870 162 19873
rect 126 19864 162 19870
rect 810 19870 816 19873
rect 810 19864 1584 19870
rect 126 19830 138 19864
rect 1572 19830 1584 19864
rect 126 19824 162 19830
rect 156 19821 162 19824
rect 810 19824 1584 19830
rect 810 19821 816 19824
rect 894 19784 900 19787
rect 126 19778 900 19784
rect 1548 19784 1554 19787
rect 1548 19778 1584 19784
rect 126 19744 138 19778
rect 1572 19744 1584 19778
rect 126 19738 900 19744
rect 894 19735 900 19738
rect 1548 19738 1584 19744
rect 1548 19735 1554 19738
rect 156 19698 162 19701
rect 126 19692 162 19698
rect 810 19698 816 19701
rect 810 19692 1584 19698
rect 126 19658 138 19692
rect 1572 19658 1584 19692
rect 126 19652 162 19658
rect 156 19649 162 19652
rect 810 19652 1584 19658
rect 810 19649 816 19652
rect 894 19612 900 19615
rect 126 19606 900 19612
rect 1548 19612 1554 19615
rect 1548 19606 1584 19612
rect 126 19572 138 19606
rect 1572 19572 1584 19606
rect 126 19566 900 19572
rect 894 19563 900 19566
rect 1548 19566 1584 19572
rect 1548 19563 1554 19566
rect 156 19526 162 19529
rect 126 19520 162 19526
rect 810 19526 816 19529
rect 810 19520 1584 19526
rect 126 19486 138 19520
rect 1572 19486 1584 19520
rect 126 19480 162 19486
rect 156 19477 162 19480
rect 810 19480 1584 19486
rect 810 19477 816 19480
rect 894 19440 900 19443
rect 126 19434 900 19440
rect 1548 19440 1554 19443
rect 1548 19434 1584 19440
rect 126 19400 138 19434
rect 1572 19400 1584 19434
rect 126 19394 900 19400
rect 894 19391 900 19394
rect 1548 19394 1584 19400
rect 1548 19391 1554 19394
rect 156 19354 162 19357
rect 126 19348 162 19354
rect 810 19354 816 19357
rect 810 19348 1584 19354
rect 126 19314 138 19348
rect 1572 19314 1584 19348
rect 126 19308 162 19314
rect 156 19305 162 19308
rect 810 19308 1584 19314
rect 810 19305 816 19308
rect 894 19268 900 19271
rect 126 19262 900 19268
rect 1548 19268 1554 19271
rect 1548 19262 1584 19268
rect 126 19228 138 19262
rect 1572 19228 1584 19262
rect 126 19222 900 19228
rect 894 19219 900 19222
rect 1548 19222 1584 19228
rect 1548 19219 1554 19222
rect 156 19182 162 19185
rect 126 19176 162 19182
rect 810 19182 816 19185
rect 810 19176 1584 19182
rect 126 19142 138 19176
rect 1572 19142 1584 19176
rect 126 19136 162 19142
rect 156 19133 162 19136
rect 810 19136 1584 19142
rect 810 19133 816 19136
rect 894 19096 900 19099
rect 126 19090 900 19096
rect 1548 19096 1554 19099
rect 1548 19090 1584 19096
rect 126 19056 138 19090
rect 1572 19056 1584 19090
rect 126 19050 900 19056
rect 894 19047 900 19050
rect 1548 19050 1584 19056
rect 1548 19047 1554 19050
rect 156 19010 162 19013
rect 126 19004 162 19010
rect 810 19010 816 19013
rect 810 19004 1584 19010
rect 126 18970 138 19004
rect 1572 18970 1584 19004
rect 126 18964 162 18970
rect 156 18961 162 18964
rect 810 18964 1584 18970
rect 810 18961 816 18964
rect 894 18924 900 18927
rect 126 18918 900 18924
rect 1548 18924 1554 18927
rect 1548 18918 1584 18924
rect 126 18884 138 18918
rect 1572 18884 1584 18918
rect 126 18878 900 18884
rect 894 18875 900 18878
rect 1548 18878 1584 18884
rect 1548 18875 1554 18878
rect 156 18838 162 18841
rect 126 18832 162 18838
rect 810 18838 816 18841
rect 810 18832 1584 18838
rect 126 18798 138 18832
rect 1572 18798 1584 18832
rect 126 18792 162 18798
rect 156 18789 162 18792
rect 810 18792 1584 18798
rect 810 18789 816 18792
rect 894 18752 900 18755
rect 126 18746 900 18752
rect 1548 18752 1554 18755
rect 1548 18746 1584 18752
rect 126 18712 138 18746
rect 1572 18712 1584 18746
rect 126 18706 900 18712
rect 894 18703 900 18706
rect 1548 18706 1584 18712
rect 1548 18703 1554 18706
rect 156 18666 162 18669
rect 126 18660 162 18666
rect 810 18666 816 18669
rect 810 18660 1584 18666
rect 126 18626 138 18660
rect 1572 18626 1584 18660
rect 126 18620 162 18626
rect 156 18617 162 18620
rect 810 18620 1584 18626
rect 810 18617 816 18620
rect 894 18580 900 18583
rect 126 18574 900 18580
rect 1548 18580 1554 18583
rect 1548 18574 1584 18580
rect 126 18540 138 18574
rect 1572 18540 1584 18574
rect 126 18534 900 18540
rect 894 18531 900 18534
rect 1548 18534 1584 18540
rect 1548 18531 1554 18534
rect 156 18494 162 18497
rect 126 18488 162 18494
rect 810 18494 816 18497
rect 810 18488 1584 18494
rect 126 18454 138 18488
rect 1572 18454 1584 18488
rect 126 18448 162 18454
rect 156 18445 162 18448
rect 810 18448 1584 18454
rect 810 18445 816 18448
rect 894 18408 900 18411
rect 126 18402 900 18408
rect 1548 18408 1554 18411
rect 1548 18402 1584 18408
rect 126 18368 138 18402
rect 1572 18368 1584 18402
rect 126 18362 900 18368
rect 894 18359 900 18362
rect 1548 18362 1584 18368
rect 1548 18359 1554 18362
rect 156 18322 162 18325
rect 126 18316 162 18322
rect 810 18322 816 18325
rect 810 18316 1584 18322
rect 126 18282 138 18316
rect 1572 18282 1584 18316
rect 126 18276 162 18282
rect 156 18273 162 18276
rect 810 18276 1584 18282
rect 810 18273 816 18276
rect 894 18236 900 18239
rect 126 18230 900 18236
rect 1548 18236 1554 18239
rect 1548 18230 1584 18236
rect 126 18196 138 18230
rect 1572 18196 1584 18230
rect 126 18190 900 18196
rect 894 18187 900 18190
rect 1548 18190 1584 18196
rect 1548 18187 1554 18190
rect 156 18150 162 18153
rect 126 18144 162 18150
rect 810 18150 816 18153
rect 810 18144 1584 18150
rect 126 18110 138 18144
rect 1572 18110 1584 18144
rect 126 18104 162 18110
rect 156 18101 162 18104
rect 810 18104 1584 18110
rect 810 18101 816 18104
rect 894 18064 900 18067
rect 126 18058 900 18064
rect 1548 18064 1554 18067
rect 1548 18058 1584 18064
rect 126 18024 138 18058
rect 1572 18024 1584 18058
rect 126 18018 900 18024
rect 894 18015 900 18018
rect 1548 18018 1584 18024
rect 1548 18015 1554 18018
rect 156 17978 162 17981
rect 126 17972 162 17978
rect 810 17978 816 17981
rect 810 17972 1584 17978
rect 126 17938 138 17972
rect 1572 17938 1584 17972
rect 126 17932 162 17938
rect 156 17929 162 17932
rect 810 17932 1584 17938
rect 810 17929 816 17932
rect 894 17892 900 17895
rect 126 17886 900 17892
rect 1548 17892 1554 17895
rect 1548 17886 1584 17892
rect 126 17852 138 17886
rect 1572 17852 1584 17886
rect 126 17846 900 17852
rect 894 17843 900 17846
rect 1548 17846 1584 17852
rect 1548 17843 1554 17846
rect 156 17806 162 17809
rect 126 17800 162 17806
rect 810 17806 816 17809
rect 810 17800 1584 17806
rect 126 17766 138 17800
rect 1572 17766 1584 17800
rect 126 17760 162 17766
rect 156 17757 162 17760
rect 810 17760 1584 17766
rect 810 17757 816 17760
rect 894 17720 900 17723
rect 126 17714 900 17720
rect 1548 17720 1554 17723
rect 1548 17714 1584 17720
rect 126 17680 138 17714
rect 1572 17680 1584 17714
rect 126 17674 900 17680
rect 894 17671 900 17674
rect 1548 17674 1584 17680
rect 1548 17671 1554 17674
rect 156 17634 162 17637
rect 126 17628 162 17634
rect 810 17634 816 17637
rect 810 17628 1584 17634
rect 126 17594 138 17628
rect 1572 17594 1584 17628
rect 126 17588 162 17594
rect 156 17585 162 17588
rect 810 17588 1584 17594
rect 810 17585 816 17588
rect 894 17548 900 17551
rect 126 17542 900 17548
rect 1548 17548 1554 17551
rect 1548 17542 1584 17548
rect 126 17508 138 17542
rect 1572 17508 1584 17542
rect 126 17502 900 17508
rect 894 17499 900 17502
rect 1548 17502 1584 17508
rect 1548 17499 1554 17502
rect 156 17462 162 17465
rect 126 17456 162 17462
rect 810 17462 816 17465
rect 810 17456 1584 17462
rect 126 17422 138 17456
rect 1572 17422 1584 17456
rect 126 17416 162 17422
rect 156 17413 162 17416
rect 810 17416 1584 17422
rect 810 17413 816 17416
rect 894 17376 900 17379
rect 126 17370 900 17376
rect 1548 17376 1554 17379
rect 1548 17370 1584 17376
rect 126 17336 138 17370
rect 1572 17336 1584 17370
rect 126 17330 900 17336
rect 894 17327 900 17330
rect 1548 17330 1584 17336
rect 1548 17327 1554 17330
rect 156 17290 162 17293
rect 126 17284 162 17290
rect 810 17290 816 17293
rect 810 17284 1584 17290
rect 126 17250 138 17284
rect 1572 17250 1584 17284
rect 126 17244 162 17250
rect 156 17241 162 17244
rect 810 17244 1584 17250
rect 810 17241 816 17244
rect 894 17204 900 17207
rect 126 17198 900 17204
rect 1548 17204 1554 17207
rect 1548 17198 1584 17204
rect 126 17164 138 17198
rect 1572 17164 1584 17198
rect 126 17158 900 17164
rect 894 17155 900 17158
rect 1548 17158 1584 17164
rect 1548 17155 1554 17158
rect 156 17118 162 17121
rect 126 17112 162 17118
rect 810 17118 816 17121
rect 810 17112 1584 17118
rect 126 17078 138 17112
rect 1572 17078 1584 17112
rect 126 17072 162 17078
rect 156 17069 162 17072
rect 810 17072 1584 17078
rect 810 17069 816 17072
rect 894 17032 900 17035
rect 126 17026 900 17032
rect 1548 17032 1554 17035
rect 1548 17026 1584 17032
rect 126 16992 138 17026
rect 1572 16992 1584 17026
rect 126 16986 900 16992
rect 894 16983 900 16986
rect 1548 16986 1584 16992
rect 1548 16983 1554 16986
rect 156 16946 162 16949
rect 126 16940 162 16946
rect 810 16946 816 16949
rect 810 16940 1584 16946
rect 126 16906 138 16940
rect 1572 16906 1584 16940
rect 126 16900 162 16906
rect 156 16897 162 16900
rect 810 16900 1584 16906
rect 810 16897 816 16900
rect 894 16860 900 16863
rect 126 16854 900 16860
rect 1548 16860 1554 16863
rect 1548 16854 1584 16860
rect 126 16820 138 16854
rect 1572 16820 1584 16854
rect 126 16814 900 16820
rect 894 16811 900 16814
rect 1548 16814 1584 16820
rect 1548 16811 1554 16814
rect 156 16774 162 16777
rect 126 16768 162 16774
rect 810 16774 816 16777
rect 810 16768 1584 16774
rect 126 16734 138 16768
rect 1572 16734 1584 16768
rect 126 16728 162 16734
rect 156 16725 162 16728
rect 810 16728 1584 16734
rect 810 16725 816 16728
rect 894 16688 900 16691
rect 126 16682 900 16688
rect 1548 16688 1554 16691
rect 1548 16682 1584 16688
rect 126 16648 138 16682
rect 1572 16648 1584 16682
rect 126 16642 900 16648
rect 894 16639 900 16642
rect 1548 16642 1584 16648
rect 1548 16639 1554 16642
rect 156 16602 162 16605
rect 126 16596 162 16602
rect 810 16602 816 16605
rect 810 16596 1584 16602
rect 126 16562 138 16596
rect 1572 16562 1584 16596
rect 126 16556 162 16562
rect 156 16553 162 16556
rect 810 16556 1584 16562
rect 810 16553 816 16556
rect 894 16516 900 16519
rect 126 16510 900 16516
rect 1548 16516 1554 16519
rect 1548 16510 1584 16516
rect 126 16476 138 16510
rect 1572 16476 1584 16510
rect 126 16470 900 16476
rect 894 16467 900 16470
rect 1548 16470 1584 16476
rect 1548 16467 1554 16470
rect 156 16430 162 16433
rect 126 16424 162 16430
rect 810 16430 816 16433
rect 810 16424 1584 16430
rect 126 16390 138 16424
rect 1572 16390 1584 16424
rect 126 16384 162 16390
rect 156 16381 162 16384
rect 810 16384 1584 16390
rect 810 16381 816 16384
rect 894 16344 900 16347
rect 126 16338 900 16344
rect 1548 16344 1554 16347
rect 1548 16338 1584 16344
rect 126 16304 138 16338
rect 1572 16304 1584 16338
rect 126 16298 900 16304
rect 894 16295 900 16298
rect 1548 16298 1584 16304
rect 1548 16295 1554 16298
rect 156 16258 162 16261
rect 126 16252 162 16258
rect 810 16258 816 16261
rect 810 16252 1584 16258
rect 126 16218 138 16252
rect 1572 16218 1584 16252
rect 126 16212 162 16218
rect 156 16209 162 16212
rect 810 16212 1584 16218
rect 810 16209 816 16212
rect 894 16172 900 16175
rect 126 16166 900 16172
rect 1548 16172 1554 16175
rect 1548 16166 1584 16172
rect 126 16132 138 16166
rect 1572 16132 1584 16166
rect 126 16126 900 16132
rect 894 16123 900 16126
rect 1548 16126 1584 16132
rect 1548 16123 1554 16126
rect 156 16086 162 16089
rect 126 16080 162 16086
rect 810 16086 816 16089
rect 810 16080 1584 16086
rect 126 16046 138 16080
rect 1572 16046 1584 16080
rect 126 16040 162 16046
rect 156 16037 162 16040
rect 810 16040 1584 16046
rect 810 16037 816 16040
rect 894 16000 900 16003
rect 126 15994 900 16000
rect 1548 16000 1554 16003
rect 1548 15994 1584 16000
rect 126 15960 138 15994
rect 1572 15960 1584 15994
rect 126 15954 900 15960
rect 894 15951 900 15954
rect 1548 15954 1584 15960
rect 1548 15951 1554 15954
rect 156 15914 162 15917
rect 126 15908 162 15914
rect 810 15914 816 15917
rect 810 15908 1584 15914
rect 126 15874 138 15908
rect 1572 15874 1584 15908
rect 126 15868 162 15874
rect 156 15865 162 15868
rect 810 15868 1584 15874
rect 810 15865 816 15868
rect 894 15828 900 15831
rect 126 15822 900 15828
rect 1548 15828 1554 15831
rect 1548 15822 1584 15828
rect 126 15788 138 15822
rect 1572 15788 1584 15822
rect 126 15782 900 15788
rect 894 15779 900 15782
rect 1548 15782 1584 15788
rect 1548 15779 1554 15782
rect 156 15742 162 15745
rect 126 15736 162 15742
rect 810 15742 816 15745
rect 810 15736 1584 15742
rect 126 15702 138 15736
rect 1572 15702 1584 15736
rect 126 15696 162 15702
rect 156 15693 162 15696
rect 810 15696 1584 15702
rect 810 15693 816 15696
rect 894 15656 900 15659
rect 126 15650 900 15656
rect 1548 15656 1554 15659
rect 1548 15650 1584 15656
rect 126 15616 138 15650
rect 1572 15616 1584 15650
rect 126 15610 900 15616
rect 894 15607 900 15610
rect 1548 15610 1584 15616
rect 1548 15607 1554 15610
rect 156 15570 162 15573
rect 126 15564 162 15570
rect 810 15570 816 15573
rect 810 15564 1584 15570
rect 126 15530 138 15564
rect 1572 15530 1584 15564
rect 126 15524 162 15530
rect 156 15521 162 15524
rect 810 15524 1584 15530
rect 810 15521 816 15524
rect 894 15484 900 15487
rect 126 15478 900 15484
rect 1548 15484 1554 15487
rect 1548 15478 1584 15484
rect 126 15444 138 15478
rect 1572 15444 1584 15478
rect 126 15438 900 15444
rect 894 15435 900 15438
rect 1548 15438 1584 15444
rect 1548 15435 1554 15438
rect 156 15398 162 15401
rect 126 15392 162 15398
rect 810 15398 816 15401
rect 810 15392 1584 15398
rect 126 15358 138 15392
rect 1572 15358 1584 15392
rect 126 15352 162 15358
rect 156 15349 162 15352
rect 810 15352 1584 15358
rect 810 15349 816 15352
rect 894 15312 900 15315
rect 126 15306 900 15312
rect 1548 15312 1554 15315
rect 1548 15306 1584 15312
rect 126 15272 138 15306
rect 1572 15272 1584 15306
rect 126 15266 900 15272
rect 894 15263 900 15266
rect 1548 15266 1584 15272
rect 1548 15263 1554 15266
rect 156 15226 162 15229
rect 126 15220 162 15226
rect 810 15226 816 15229
rect 810 15220 1584 15226
rect 126 15186 138 15220
rect 1572 15186 1584 15220
rect 126 15180 162 15186
rect 156 15177 162 15180
rect 810 15180 1584 15186
rect 810 15177 816 15180
rect 894 15140 900 15143
rect 126 15134 900 15140
rect 1548 15140 1554 15143
rect 1548 15134 1584 15140
rect 126 15100 138 15134
rect 1572 15100 1584 15134
rect 126 15094 900 15100
rect 894 15091 900 15094
rect 1548 15094 1584 15100
rect 1548 15091 1554 15094
rect 156 15054 162 15057
rect 126 15048 162 15054
rect 810 15054 816 15057
rect 810 15048 1584 15054
rect 126 15014 138 15048
rect 1572 15014 1584 15048
rect 126 15008 162 15014
rect 156 15005 162 15008
rect 810 15008 1584 15014
rect 810 15005 816 15008
rect 894 14968 900 14971
rect 126 14962 900 14968
rect 1548 14968 1554 14971
rect 1548 14962 1584 14968
rect 126 14928 138 14962
rect 1572 14928 1584 14962
rect 126 14922 900 14928
rect 894 14919 900 14922
rect 1548 14922 1584 14928
rect 1548 14919 1554 14922
rect 156 14882 162 14885
rect 126 14876 162 14882
rect 810 14882 816 14885
rect 810 14876 1584 14882
rect 126 14842 138 14876
rect 1572 14842 1584 14876
rect 126 14836 162 14842
rect 156 14833 162 14836
rect 810 14836 1584 14842
rect 810 14833 816 14836
rect 894 14796 900 14799
rect 126 14790 900 14796
rect 1548 14796 1554 14799
rect 1548 14790 1584 14796
rect 126 14756 138 14790
rect 1572 14756 1584 14790
rect 126 14750 900 14756
rect 894 14747 900 14750
rect 1548 14750 1584 14756
rect 1548 14747 1554 14750
rect 156 14710 162 14713
rect 126 14704 162 14710
rect 810 14710 816 14713
rect 810 14704 1584 14710
rect 126 14670 138 14704
rect 1572 14670 1584 14704
rect 126 14664 162 14670
rect 156 14661 162 14664
rect 810 14664 1584 14670
rect 810 14661 816 14664
rect 894 14624 900 14627
rect 126 14618 900 14624
rect 1548 14624 1554 14627
rect 1548 14618 1584 14624
rect 126 14584 138 14618
rect 1572 14584 1584 14618
rect 126 14578 900 14584
rect 894 14575 900 14578
rect 1548 14578 1584 14584
rect 1548 14575 1554 14578
rect 156 14538 162 14541
rect 126 14532 162 14538
rect 810 14538 816 14541
rect 810 14532 1584 14538
rect 126 14498 138 14532
rect 1572 14498 1584 14532
rect 126 14492 162 14498
rect 156 14489 162 14492
rect 810 14492 1584 14498
rect 810 14489 816 14492
rect 894 14452 900 14455
rect 126 14446 900 14452
rect 1548 14452 1554 14455
rect 1548 14446 1584 14452
rect 126 14412 138 14446
rect 1572 14412 1584 14446
rect 126 14406 900 14412
rect 894 14403 900 14406
rect 1548 14406 1584 14412
rect 1548 14403 1554 14406
rect 156 14366 162 14369
rect 126 14360 162 14366
rect 810 14366 816 14369
rect 810 14360 1584 14366
rect 126 14326 138 14360
rect 1572 14326 1584 14360
rect 126 14320 162 14326
rect 156 14317 162 14320
rect 810 14320 1584 14326
rect 810 14317 816 14320
rect 894 14280 900 14283
rect 126 14274 900 14280
rect 1548 14280 1554 14283
rect 1548 14274 1584 14280
rect 126 14240 138 14274
rect 1572 14240 1584 14274
rect 126 14234 900 14240
rect 894 14231 900 14234
rect 1548 14234 1584 14240
rect 1548 14231 1554 14234
rect 156 14194 162 14197
rect 126 14188 162 14194
rect 810 14194 816 14197
rect 810 14188 1584 14194
rect 126 14154 138 14188
rect 1572 14154 1584 14188
rect 126 14148 162 14154
rect 156 14145 162 14148
rect 810 14148 1584 14154
rect 810 14145 816 14148
rect 894 14108 900 14111
rect 126 14102 900 14108
rect 1548 14108 1554 14111
rect 1548 14102 1584 14108
rect 126 14068 138 14102
rect 1572 14068 1584 14102
rect 126 14062 900 14068
rect 894 14059 900 14062
rect 1548 14062 1584 14068
rect 1548 14059 1554 14062
rect 156 14022 162 14025
rect 126 14016 162 14022
rect 810 14022 816 14025
rect 810 14016 1584 14022
rect 126 13982 138 14016
rect 1572 13982 1584 14016
rect 126 13976 162 13982
rect 156 13973 162 13976
rect 810 13976 1584 13982
rect 810 13973 816 13976
rect 894 13936 900 13939
rect 126 13930 900 13936
rect 1548 13936 1554 13939
rect 1548 13930 1584 13936
rect 126 13896 138 13930
rect 1572 13896 1584 13930
rect 126 13890 900 13896
rect 894 13887 900 13890
rect 1548 13890 1584 13896
rect 1548 13887 1554 13890
rect 156 13850 162 13853
rect 126 13844 162 13850
rect 810 13850 816 13853
rect 810 13844 1584 13850
rect 126 13810 138 13844
rect 1572 13810 1584 13844
rect 126 13804 162 13810
rect 156 13801 162 13804
rect 810 13804 1584 13810
rect 810 13801 816 13804
rect 894 13764 900 13767
rect 126 13758 900 13764
rect 1548 13764 1554 13767
rect 1548 13758 1584 13764
rect 126 13724 138 13758
rect 1572 13724 1584 13758
rect 126 13718 900 13724
rect 894 13715 900 13718
rect 1548 13718 1584 13724
rect 1548 13715 1554 13718
rect 156 13678 162 13681
rect 126 13672 162 13678
rect 810 13678 816 13681
rect 810 13672 1584 13678
rect 126 13638 138 13672
rect 1572 13638 1584 13672
rect 126 13632 162 13638
rect 156 13629 162 13632
rect 810 13632 1584 13638
rect 810 13629 816 13632
rect 894 13592 900 13595
rect 126 13586 900 13592
rect 1548 13592 1554 13595
rect 1548 13586 1584 13592
rect 126 13552 138 13586
rect 1572 13552 1584 13586
rect 126 13546 900 13552
rect 894 13543 900 13546
rect 1548 13546 1584 13552
rect 1548 13543 1554 13546
rect 156 13506 162 13509
rect 126 13500 162 13506
rect 810 13506 816 13509
rect 810 13500 1584 13506
rect 126 13466 138 13500
rect 1572 13466 1584 13500
rect 126 13460 162 13466
rect 156 13457 162 13460
rect 810 13460 1584 13466
rect 810 13457 816 13460
rect 894 13420 900 13423
rect 126 13414 900 13420
rect 1548 13420 1554 13423
rect 1548 13414 1584 13420
rect 126 13380 138 13414
rect 1572 13380 1584 13414
rect 126 13374 900 13380
rect 894 13371 900 13374
rect 1548 13374 1584 13380
rect 1548 13371 1554 13374
rect 156 13334 162 13337
rect 126 13328 162 13334
rect 810 13334 816 13337
rect 810 13328 1584 13334
rect 126 13294 138 13328
rect 1572 13294 1584 13328
rect 126 13288 162 13294
rect 156 13285 162 13288
rect 810 13288 1584 13294
rect 810 13285 816 13288
rect 894 13248 900 13251
rect 126 13242 900 13248
rect 1548 13248 1554 13251
rect 1548 13242 1584 13248
rect 126 13208 138 13242
rect 1572 13208 1584 13242
rect 126 13202 900 13208
rect 894 13199 900 13202
rect 1548 13202 1584 13208
rect 1548 13199 1554 13202
rect 156 13162 162 13165
rect 126 13156 162 13162
rect 810 13162 816 13165
rect 810 13156 1584 13162
rect 126 13122 138 13156
rect 1572 13122 1584 13156
rect 126 13116 162 13122
rect 156 13113 162 13116
rect 810 13116 1584 13122
rect 810 13113 816 13116
rect 894 13076 900 13079
rect 126 13070 900 13076
rect 1548 13076 1554 13079
rect 1548 13070 1584 13076
rect 126 13036 138 13070
rect 1572 13036 1584 13070
rect 126 13030 900 13036
rect 894 13027 900 13030
rect 1548 13030 1584 13036
rect 1548 13027 1554 13030
rect 156 12990 162 12993
rect 126 12984 162 12990
rect 810 12990 816 12993
rect 810 12984 1584 12990
rect 126 12950 138 12984
rect 1572 12950 1584 12984
rect 126 12944 162 12950
rect 156 12941 162 12944
rect 810 12944 1584 12950
rect 810 12941 816 12944
rect 894 12904 900 12907
rect 126 12898 900 12904
rect 1548 12904 1554 12907
rect 1548 12898 1584 12904
rect 126 12864 138 12898
rect 1572 12864 1584 12898
rect 126 12858 900 12864
rect 894 12855 900 12858
rect 1548 12858 1584 12864
rect 1548 12855 1554 12858
rect 156 12818 162 12821
rect 126 12812 162 12818
rect 810 12818 816 12821
rect 810 12812 1584 12818
rect 126 12778 138 12812
rect 1572 12778 1584 12812
rect 126 12772 162 12778
rect 156 12769 162 12772
rect 810 12772 1584 12778
rect 810 12769 816 12772
rect 894 12732 900 12735
rect 126 12726 900 12732
rect 1548 12732 1554 12735
rect 1548 12726 1584 12732
rect 126 12692 138 12726
rect 1572 12692 1584 12726
rect 126 12686 900 12692
rect 894 12683 900 12686
rect 1548 12686 1584 12692
rect 1548 12683 1554 12686
rect 156 12646 162 12649
rect 126 12640 162 12646
rect 810 12646 816 12649
rect 810 12640 1584 12646
rect 126 12606 138 12640
rect 1572 12606 1584 12640
rect 126 12600 162 12606
rect 156 12597 162 12600
rect 810 12600 1584 12606
rect 810 12597 816 12600
rect 894 12560 900 12563
rect 126 12554 900 12560
rect 1548 12560 1554 12563
rect 1548 12554 1584 12560
rect 126 12520 138 12554
rect 1572 12520 1584 12554
rect 126 12514 900 12520
rect 894 12511 900 12514
rect 1548 12514 1584 12520
rect 1548 12511 1554 12514
rect 156 12474 162 12477
rect 126 12468 162 12474
rect 810 12474 816 12477
rect 810 12468 1584 12474
rect 126 12434 138 12468
rect 1572 12434 1584 12468
rect 126 12428 162 12434
rect 156 12425 162 12428
rect 810 12428 1584 12434
rect 810 12425 816 12428
rect 894 12388 900 12391
rect 126 12382 900 12388
rect 1548 12388 1554 12391
rect 1548 12382 1584 12388
rect 126 12348 138 12382
rect 1572 12348 1584 12382
rect 126 12342 900 12348
rect 894 12339 900 12342
rect 1548 12342 1584 12348
rect 1548 12339 1554 12342
rect 156 12302 162 12305
rect 126 12296 162 12302
rect 810 12302 816 12305
rect 810 12296 1584 12302
rect 126 12262 138 12296
rect 1572 12262 1584 12296
rect 126 12256 162 12262
rect 156 12253 162 12256
rect 810 12256 1584 12262
rect 810 12253 816 12256
rect 894 12216 900 12219
rect 126 12210 900 12216
rect 1548 12216 1554 12219
rect 1548 12210 1584 12216
rect 126 12176 138 12210
rect 1572 12176 1584 12210
rect 126 12170 900 12176
rect 894 12167 900 12170
rect 1548 12170 1584 12176
rect 1548 12167 1554 12170
rect 156 12130 162 12133
rect 126 12124 162 12130
rect 810 12130 816 12133
rect 810 12124 1584 12130
rect 126 12090 138 12124
rect 1572 12090 1584 12124
rect 126 12084 162 12090
rect 156 12081 162 12084
rect 810 12084 1584 12090
rect 810 12081 816 12084
rect 894 12044 900 12047
rect 126 12038 900 12044
rect 1548 12044 1554 12047
rect 1548 12038 1584 12044
rect 126 12004 138 12038
rect 1572 12004 1584 12038
rect 126 11998 900 12004
rect 894 11995 900 11998
rect 1548 11998 1584 12004
rect 1548 11995 1554 11998
rect 156 11958 162 11961
rect 126 11952 162 11958
rect 810 11958 816 11961
rect 810 11952 1584 11958
rect 126 11918 138 11952
rect 1572 11918 1584 11952
rect 126 11912 162 11918
rect 156 11909 162 11912
rect 810 11912 1584 11918
rect 810 11909 816 11912
rect 894 11872 900 11875
rect 126 11866 900 11872
rect 1548 11872 1554 11875
rect 1548 11866 1584 11872
rect 126 11832 138 11866
rect 1572 11832 1584 11866
rect 126 11826 900 11832
rect 894 11823 900 11826
rect 1548 11826 1584 11832
rect 1548 11823 1554 11826
rect 156 11786 162 11789
rect 126 11780 162 11786
rect 810 11786 816 11789
rect 810 11780 1584 11786
rect 126 11746 138 11780
rect 1572 11746 1584 11780
rect 126 11740 162 11746
rect 156 11737 162 11740
rect 810 11740 1584 11746
rect 810 11737 816 11740
rect 894 11700 900 11703
rect 126 11694 900 11700
rect 1548 11700 1554 11703
rect 1548 11694 1584 11700
rect 126 11660 138 11694
rect 1572 11660 1584 11694
rect 126 11654 900 11660
rect 894 11651 900 11654
rect 1548 11654 1584 11660
rect 1548 11651 1554 11654
rect 156 11614 162 11617
rect 126 11608 162 11614
rect 810 11614 816 11617
rect 810 11608 1584 11614
rect 126 11574 138 11608
rect 1572 11574 1584 11608
rect 126 11568 162 11574
rect 156 11565 162 11568
rect 810 11568 1584 11574
rect 810 11565 816 11568
rect 894 11528 900 11531
rect 126 11522 900 11528
rect 1548 11528 1554 11531
rect 1548 11522 1584 11528
rect 126 11488 138 11522
rect 1572 11488 1584 11522
rect 126 11482 900 11488
rect 894 11479 900 11482
rect 1548 11482 1584 11488
rect 1548 11479 1554 11482
rect 156 11442 162 11445
rect 126 11436 162 11442
rect 810 11442 816 11445
rect 810 11436 1584 11442
rect 126 11402 138 11436
rect 1572 11402 1584 11436
rect 126 11396 162 11402
rect 156 11393 162 11396
rect 810 11396 1584 11402
rect 810 11393 816 11396
rect 894 11356 900 11359
rect 126 11350 900 11356
rect 1548 11356 1554 11359
rect 1548 11350 1584 11356
rect 126 11316 138 11350
rect 1572 11316 1584 11350
rect 126 11310 900 11316
rect 894 11307 900 11310
rect 1548 11310 1584 11316
rect 1548 11307 1554 11310
rect 156 11270 162 11273
rect 126 11264 162 11270
rect 810 11270 816 11273
rect 810 11264 1584 11270
rect 126 11230 138 11264
rect 1572 11230 1584 11264
rect 126 11224 162 11230
rect 156 11221 162 11224
rect 810 11224 1584 11230
rect 810 11221 816 11224
rect 894 11184 900 11187
rect 126 11178 900 11184
rect 1548 11184 1554 11187
rect 1548 11178 1584 11184
rect 126 11144 138 11178
rect 1572 11144 1584 11178
rect 126 11138 900 11144
rect 894 11135 900 11138
rect 1548 11138 1584 11144
rect 1548 11135 1554 11138
rect 156 11098 162 11101
rect 126 11092 162 11098
rect 810 11098 816 11101
rect 810 11092 1584 11098
rect 126 11058 138 11092
rect 1572 11058 1584 11092
rect 126 11052 162 11058
rect 156 11049 162 11052
rect 810 11052 1584 11058
rect 810 11049 816 11052
rect 894 11012 900 11015
rect 126 11006 900 11012
rect 1548 11012 1554 11015
rect 1548 11006 1584 11012
rect 126 10972 138 11006
rect 1572 10972 1584 11006
rect 126 10966 900 10972
rect 894 10963 900 10966
rect 1548 10966 1584 10972
rect 1548 10963 1554 10966
rect 156 10926 162 10929
rect 126 10920 162 10926
rect 810 10926 816 10929
rect 810 10920 1584 10926
rect 126 10886 138 10920
rect 1572 10886 1584 10920
rect 126 10880 162 10886
rect 156 10877 162 10880
rect 810 10880 1584 10886
rect 810 10877 816 10880
rect 894 10840 900 10843
rect 126 10834 900 10840
rect 1548 10840 1554 10843
rect 1548 10834 1584 10840
rect 126 10800 138 10834
rect 1572 10800 1584 10834
rect 126 10794 900 10800
rect 894 10791 900 10794
rect 1548 10794 1584 10800
rect 1548 10791 1554 10794
rect 156 10754 162 10757
rect 126 10748 162 10754
rect 810 10754 816 10757
rect 810 10748 1584 10754
rect 126 10714 138 10748
rect 1572 10714 1584 10748
rect 126 10708 162 10714
rect 156 10705 162 10708
rect 810 10708 1584 10714
rect 810 10705 816 10708
rect 894 10668 900 10671
rect 126 10662 900 10668
rect 1548 10668 1554 10671
rect 1548 10662 1584 10668
rect 126 10628 138 10662
rect 1572 10628 1584 10662
rect 126 10622 900 10628
rect 894 10619 900 10622
rect 1548 10622 1584 10628
rect 1548 10619 1554 10622
rect 156 10582 162 10585
rect 126 10576 162 10582
rect 810 10582 816 10585
rect 810 10576 1584 10582
rect 126 10542 138 10576
rect 1572 10542 1584 10576
rect 126 10536 162 10542
rect 156 10533 162 10536
rect 810 10536 1584 10542
rect 810 10533 816 10536
rect 894 10496 900 10499
rect 126 10490 900 10496
rect 1548 10496 1554 10499
rect 1548 10490 1584 10496
rect 126 10456 138 10490
rect 1572 10456 1584 10490
rect 126 10450 900 10456
rect 894 10447 900 10450
rect 1548 10450 1584 10456
rect 1548 10447 1554 10450
rect 156 10410 162 10413
rect 126 10404 162 10410
rect 810 10410 816 10413
rect 810 10404 1584 10410
rect 126 10370 138 10404
rect 1572 10370 1584 10404
rect 126 10364 162 10370
rect 156 10361 162 10364
rect 810 10364 1584 10370
rect 810 10361 816 10364
rect 894 10324 900 10327
rect 126 10318 900 10324
rect 1548 10324 1554 10327
rect 1548 10318 1584 10324
rect 126 10284 138 10318
rect 1572 10284 1584 10318
rect 126 10278 900 10284
rect 894 10275 900 10278
rect 1548 10278 1584 10284
rect 1548 10275 1554 10278
rect 156 10238 162 10241
rect 126 10232 162 10238
rect 810 10238 816 10241
rect 810 10232 1584 10238
rect 126 10198 138 10232
rect 1572 10198 1584 10232
rect 126 10192 162 10198
rect 156 10189 162 10192
rect 810 10192 1584 10198
rect 810 10189 816 10192
rect 894 10152 900 10155
rect 126 10146 900 10152
rect 1548 10152 1554 10155
rect 1548 10146 1584 10152
rect 126 10112 138 10146
rect 1572 10112 1584 10146
rect 126 10106 900 10112
rect 894 10103 900 10106
rect 1548 10106 1584 10112
rect 1548 10103 1554 10106
rect 156 10066 162 10069
rect 126 10060 162 10066
rect 810 10066 816 10069
rect 810 10060 1584 10066
rect 126 10026 138 10060
rect 1572 10026 1584 10060
rect 126 10020 162 10026
rect 156 10017 162 10020
rect 810 10020 1584 10026
rect 810 10017 816 10020
rect 894 9980 900 9983
rect 126 9974 900 9980
rect 1548 9980 1554 9983
rect 1548 9974 1584 9980
rect 126 9940 138 9974
rect 1572 9940 1584 9974
rect 126 9934 900 9940
rect 894 9931 900 9934
rect 1548 9934 1584 9940
rect 1548 9931 1554 9934
rect 156 9894 162 9897
rect 126 9888 162 9894
rect 810 9894 816 9897
rect 810 9888 1584 9894
rect 126 9854 138 9888
rect 1572 9854 1584 9888
rect 126 9848 162 9854
rect 156 9845 162 9848
rect 810 9848 1584 9854
rect 810 9845 816 9848
rect 894 9808 900 9811
rect 126 9802 900 9808
rect 1548 9808 1554 9811
rect 1548 9802 1584 9808
rect 126 9768 138 9802
rect 1572 9768 1584 9802
rect 126 9762 900 9768
rect 894 9759 900 9762
rect 1548 9762 1584 9768
rect 1548 9759 1554 9762
rect 156 9722 162 9725
rect 126 9716 162 9722
rect 810 9722 816 9725
rect 810 9716 1584 9722
rect 126 9682 138 9716
rect 1572 9682 1584 9716
rect 126 9676 162 9682
rect 156 9673 162 9676
rect 810 9676 1584 9682
rect 810 9673 816 9676
rect 894 9636 900 9639
rect 126 9630 900 9636
rect 1548 9636 1554 9639
rect 1548 9630 1584 9636
rect 126 9596 138 9630
rect 1572 9596 1584 9630
rect 126 9590 900 9596
rect 894 9587 900 9590
rect 1548 9590 1584 9596
rect 1548 9587 1554 9590
rect 156 9550 162 9553
rect 126 9544 162 9550
rect 810 9550 816 9553
rect 810 9544 1584 9550
rect 126 9510 138 9544
rect 1572 9510 1584 9544
rect 126 9504 162 9510
rect 156 9501 162 9504
rect 810 9504 1584 9510
rect 810 9501 816 9504
rect 894 9464 900 9467
rect 126 9458 900 9464
rect 1548 9464 1554 9467
rect 1548 9458 1584 9464
rect 126 9424 138 9458
rect 1572 9424 1584 9458
rect 126 9418 900 9424
rect 894 9415 900 9418
rect 1548 9418 1584 9424
rect 1548 9415 1554 9418
rect 156 9378 162 9381
rect 126 9372 162 9378
rect 810 9378 816 9381
rect 810 9372 1584 9378
rect 126 9338 138 9372
rect 1572 9338 1584 9372
rect 126 9332 162 9338
rect 156 9329 162 9332
rect 810 9332 1584 9338
rect 810 9329 816 9332
rect 894 9292 900 9295
rect 126 9286 900 9292
rect 1548 9292 1554 9295
rect 1548 9286 1584 9292
rect 126 9252 138 9286
rect 1572 9252 1584 9286
rect 126 9246 900 9252
rect 894 9243 900 9246
rect 1548 9246 1584 9252
rect 1548 9243 1554 9246
rect 156 9206 162 9209
rect 126 9200 162 9206
rect 810 9206 816 9209
rect 810 9200 1584 9206
rect 126 9166 138 9200
rect 1572 9166 1584 9200
rect 126 9160 162 9166
rect 156 9157 162 9160
rect 810 9160 1584 9166
rect 810 9157 816 9160
rect 894 9120 900 9123
rect 126 9114 900 9120
rect 1548 9120 1554 9123
rect 1548 9114 1584 9120
rect 126 9080 138 9114
rect 1572 9080 1584 9114
rect 126 9074 900 9080
rect 894 9071 900 9074
rect 1548 9074 1584 9080
rect 1548 9071 1554 9074
rect 156 9034 162 9037
rect 126 9028 162 9034
rect 810 9034 816 9037
rect 810 9028 1584 9034
rect 126 8994 138 9028
rect 1572 8994 1584 9028
rect 126 8988 162 8994
rect 156 8985 162 8988
rect 810 8988 1584 8994
rect 810 8985 816 8988
rect 894 8948 900 8951
rect 126 8942 900 8948
rect 1548 8948 1554 8951
rect 1548 8942 1584 8948
rect 126 8908 138 8942
rect 1572 8908 1584 8942
rect 126 8902 900 8908
rect 894 8899 900 8902
rect 1548 8902 1584 8908
rect 1548 8899 1554 8902
rect 156 8862 162 8865
rect 126 8856 162 8862
rect 810 8862 816 8865
rect 810 8856 1584 8862
rect 126 8822 138 8856
rect 1572 8822 1584 8856
rect 126 8816 162 8822
rect 156 8813 162 8816
rect 810 8816 1584 8822
rect 810 8813 816 8816
rect 894 8776 900 8779
rect 126 8770 900 8776
rect 1548 8776 1554 8779
rect 1548 8770 1584 8776
rect 126 8736 138 8770
rect 1572 8736 1584 8770
rect 126 8730 900 8736
rect 894 8727 900 8730
rect 1548 8730 1584 8736
rect 1548 8727 1554 8730
rect 156 8690 162 8693
rect 126 8684 162 8690
rect 810 8690 816 8693
rect 810 8684 1584 8690
rect 126 8650 138 8684
rect 1572 8650 1584 8684
rect 126 8644 162 8650
rect 156 8641 162 8644
rect 810 8644 1584 8650
rect 810 8641 816 8644
rect 894 8604 900 8607
rect 126 8598 900 8604
rect 1548 8604 1554 8607
rect 1548 8598 1584 8604
rect 126 8564 138 8598
rect 1572 8564 1584 8598
rect 126 8558 900 8564
rect 894 8555 900 8558
rect 1548 8558 1584 8564
rect 1548 8555 1554 8558
rect 156 8518 162 8521
rect 126 8512 162 8518
rect 810 8518 816 8521
rect 810 8512 1584 8518
rect 126 8478 138 8512
rect 1572 8478 1584 8512
rect 126 8472 162 8478
rect 156 8469 162 8472
rect 810 8472 1584 8478
rect 810 8469 816 8472
rect 894 8432 900 8435
rect 126 8426 900 8432
rect 1548 8432 1554 8435
rect 1548 8426 1584 8432
rect 126 8392 138 8426
rect 1572 8392 1584 8426
rect 126 8386 900 8392
rect 894 8383 900 8386
rect 1548 8386 1584 8392
rect 1548 8383 1554 8386
rect 156 8346 162 8349
rect 126 8340 162 8346
rect 810 8346 816 8349
rect 810 8340 1584 8346
rect 126 8306 138 8340
rect 1572 8306 1584 8340
rect 126 8300 162 8306
rect 156 8297 162 8300
rect 810 8300 1584 8306
rect 810 8297 816 8300
rect 894 8260 900 8263
rect 126 8254 900 8260
rect 1548 8260 1554 8263
rect 1548 8254 1584 8260
rect 126 8220 138 8254
rect 1572 8220 1584 8254
rect 126 8214 900 8220
rect 894 8211 900 8214
rect 1548 8214 1584 8220
rect 1548 8211 1554 8214
rect 156 8174 162 8177
rect 126 8168 162 8174
rect 810 8174 816 8177
rect 810 8168 1584 8174
rect 126 8134 138 8168
rect 1572 8134 1584 8168
rect 126 8128 162 8134
rect 156 8125 162 8128
rect 810 8128 1584 8134
rect 810 8125 816 8128
rect 894 8088 900 8091
rect 126 8082 900 8088
rect 1548 8088 1554 8091
rect 1548 8082 1584 8088
rect 126 8048 138 8082
rect 1572 8048 1584 8082
rect 126 8042 900 8048
rect 894 8039 900 8042
rect 1548 8042 1584 8048
rect 1548 8039 1554 8042
rect 156 8002 162 8005
rect 126 7996 162 8002
rect 810 8002 816 8005
rect 810 7996 1584 8002
rect 126 7962 138 7996
rect 1572 7962 1584 7996
rect 126 7956 162 7962
rect 156 7953 162 7956
rect 810 7956 1584 7962
rect 810 7953 816 7956
rect 894 7916 900 7919
rect 126 7910 900 7916
rect 1548 7916 1554 7919
rect 1548 7910 1584 7916
rect 126 7876 138 7910
rect 1572 7876 1584 7910
rect 126 7870 900 7876
rect 894 7867 900 7870
rect 1548 7870 1584 7876
rect 1548 7867 1554 7870
rect 156 7830 162 7833
rect 126 7824 162 7830
rect 810 7830 816 7833
rect 810 7824 1584 7830
rect 126 7790 138 7824
rect 1572 7790 1584 7824
rect 126 7784 162 7790
rect 156 7781 162 7784
rect 810 7784 1584 7790
rect 810 7781 816 7784
rect 894 7744 900 7747
rect 126 7738 900 7744
rect 1548 7744 1554 7747
rect 1548 7738 1584 7744
rect 126 7704 138 7738
rect 1572 7704 1584 7738
rect 126 7698 900 7704
rect 894 7695 900 7698
rect 1548 7698 1584 7704
rect 1548 7695 1554 7698
rect 156 7658 162 7661
rect 126 7652 162 7658
rect 810 7658 816 7661
rect 810 7652 1584 7658
rect 126 7618 138 7652
rect 1572 7618 1584 7652
rect 126 7612 162 7618
rect 156 7609 162 7612
rect 810 7612 1584 7618
rect 810 7609 816 7612
rect 894 7572 900 7575
rect 126 7566 900 7572
rect 1548 7572 1554 7575
rect 1548 7566 1584 7572
rect 126 7532 138 7566
rect 1572 7532 1584 7566
rect 126 7526 900 7532
rect 894 7523 900 7526
rect 1548 7526 1584 7532
rect 1548 7523 1554 7526
rect 156 7486 162 7489
rect 126 7480 162 7486
rect 810 7486 816 7489
rect 810 7480 1584 7486
rect 126 7446 138 7480
rect 1572 7446 1584 7480
rect 126 7440 162 7446
rect 156 7437 162 7440
rect 810 7440 1584 7446
rect 810 7437 816 7440
rect 894 7400 900 7403
rect 126 7394 900 7400
rect 1548 7400 1554 7403
rect 1548 7394 1584 7400
rect 126 7360 138 7394
rect 1572 7360 1584 7394
rect 126 7354 900 7360
rect 894 7351 900 7354
rect 1548 7354 1584 7360
rect 1548 7351 1554 7354
rect 156 7314 162 7317
rect 126 7308 162 7314
rect 810 7314 816 7317
rect 810 7308 1584 7314
rect 126 7274 138 7308
rect 1572 7274 1584 7308
rect 126 7268 162 7274
rect 156 7265 162 7268
rect 810 7268 1584 7274
rect 810 7265 816 7268
rect 894 7228 900 7231
rect 126 7222 900 7228
rect 1548 7228 1554 7231
rect 1548 7222 1584 7228
rect 126 7188 138 7222
rect 1572 7188 1584 7222
rect 126 7182 900 7188
rect 894 7179 900 7182
rect 1548 7182 1584 7188
rect 1548 7179 1554 7182
rect 156 7142 162 7145
rect 126 7136 162 7142
rect 810 7142 816 7145
rect 810 7136 1584 7142
rect 126 7102 138 7136
rect 1572 7102 1584 7136
rect 126 7096 162 7102
rect 156 7093 162 7096
rect 810 7096 1584 7102
rect 810 7093 816 7096
rect 894 7056 900 7059
rect 126 7050 900 7056
rect 1548 7056 1554 7059
rect 1548 7050 1584 7056
rect 126 7016 138 7050
rect 1572 7016 1584 7050
rect 126 7010 900 7016
rect 894 7007 900 7010
rect 1548 7010 1584 7016
rect 1548 7007 1554 7010
rect 156 6970 162 6973
rect 126 6964 162 6970
rect 810 6970 816 6973
rect 810 6964 1584 6970
rect 126 6930 138 6964
rect 1572 6930 1584 6964
rect 126 6924 162 6930
rect 156 6921 162 6924
rect 810 6924 1584 6930
rect 810 6921 816 6924
rect 894 6884 900 6887
rect 126 6878 900 6884
rect 1548 6884 1554 6887
rect 1548 6878 1584 6884
rect 126 6844 138 6878
rect 1572 6844 1584 6878
rect 126 6838 900 6844
rect 894 6835 900 6838
rect 1548 6838 1584 6844
rect 1548 6835 1554 6838
rect 156 6798 162 6801
rect 126 6792 162 6798
rect 810 6798 816 6801
rect 810 6792 1584 6798
rect 126 6758 138 6792
rect 1572 6758 1584 6792
rect 126 6752 162 6758
rect 156 6749 162 6752
rect 810 6752 1584 6758
rect 810 6749 816 6752
rect 894 6712 900 6715
rect 126 6706 900 6712
rect 1548 6712 1554 6715
rect 1548 6706 1584 6712
rect 126 6672 138 6706
rect 1572 6672 1584 6706
rect 126 6666 900 6672
rect 894 6663 900 6666
rect 1548 6666 1584 6672
rect 1548 6663 1554 6666
rect 156 6626 162 6629
rect 126 6620 162 6626
rect 810 6626 816 6629
rect 810 6620 1584 6626
rect 126 6586 138 6620
rect 1572 6586 1584 6620
rect 126 6580 162 6586
rect 156 6577 162 6580
rect 810 6580 1584 6586
rect 810 6577 816 6580
rect 894 6540 900 6543
rect 126 6534 900 6540
rect 1548 6540 1554 6543
rect 1548 6534 1584 6540
rect 126 6500 138 6534
rect 1572 6500 1584 6534
rect 126 6494 900 6500
rect 894 6491 900 6494
rect 1548 6494 1584 6500
rect 1548 6491 1554 6494
rect 156 6454 162 6457
rect 126 6448 162 6454
rect 810 6454 816 6457
rect 810 6448 1584 6454
rect 126 6414 138 6448
rect 1572 6414 1584 6448
rect 126 6408 162 6414
rect 156 6405 162 6408
rect 810 6408 1584 6414
rect 810 6405 816 6408
rect 894 6368 900 6371
rect 126 6362 900 6368
rect 1548 6368 1554 6371
rect 1548 6362 1584 6368
rect 126 6328 138 6362
rect 1572 6328 1584 6362
rect 126 6322 900 6328
rect 894 6319 900 6322
rect 1548 6322 1584 6328
rect 1548 6319 1554 6322
rect 156 6282 162 6285
rect 126 6276 162 6282
rect 810 6282 816 6285
rect 810 6276 1584 6282
rect 126 6242 138 6276
rect 1572 6242 1584 6276
rect 126 6236 162 6242
rect 156 6233 162 6236
rect 810 6236 1584 6242
rect 810 6233 816 6236
rect 894 6196 900 6199
rect 126 6190 900 6196
rect 1548 6196 1554 6199
rect 1548 6190 1584 6196
rect 126 6156 138 6190
rect 1572 6156 1584 6190
rect 126 6150 900 6156
rect 894 6147 900 6150
rect 1548 6150 1584 6156
rect 1548 6147 1554 6150
rect 156 6110 162 6113
rect 126 6104 162 6110
rect 810 6110 816 6113
rect 810 6104 1584 6110
rect 126 6070 138 6104
rect 1572 6070 1584 6104
rect 126 6064 162 6070
rect 156 6061 162 6064
rect 810 6064 1584 6070
rect 810 6061 816 6064
rect 894 6024 900 6027
rect 126 6018 900 6024
rect 1548 6024 1554 6027
rect 1548 6018 1584 6024
rect 126 5984 138 6018
rect 1572 5984 1584 6018
rect 126 5978 900 5984
rect 894 5975 900 5978
rect 1548 5978 1584 5984
rect 1548 5975 1554 5978
rect 156 5938 162 5941
rect 126 5932 162 5938
rect 810 5938 816 5941
rect 810 5932 1584 5938
rect 126 5898 138 5932
rect 1572 5898 1584 5932
rect 126 5892 162 5898
rect 156 5889 162 5892
rect 810 5892 1584 5898
rect 810 5889 816 5892
rect 894 5852 900 5855
rect 126 5846 900 5852
rect 1548 5852 1554 5855
rect 1548 5846 1584 5852
rect 126 5812 138 5846
rect 1572 5812 1584 5846
rect 126 5806 900 5812
rect 894 5803 900 5806
rect 1548 5806 1584 5812
rect 1548 5803 1554 5806
rect 156 5766 162 5769
rect 126 5760 162 5766
rect 810 5766 816 5769
rect 810 5760 1584 5766
rect 126 5726 138 5760
rect 1572 5726 1584 5760
rect 126 5720 162 5726
rect 156 5717 162 5720
rect 810 5720 1584 5726
rect 810 5717 816 5720
rect 894 5680 900 5683
rect 126 5674 900 5680
rect 1548 5680 1554 5683
rect 1548 5674 1584 5680
rect 126 5640 138 5674
rect 1572 5640 1584 5674
rect 126 5634 900 5640
rect 894 5631 900 5634
rect 1548 5634 1584 5640
rect 1548 5631 1554 5634
rect 156 5594 162 5597
rect 126 5588 162 5594
rect 810 5594 816 5597
rect 810 5588 1584 5594
rect 126 5554 138 5588
rect 1572 5554 1584 5588
rect 126 5548 162 5554
rect 156 5545 162 5548
rect 810 5548 1584 5554
rect 810 5545 816 5548
rect 894 5508 900 5511
rect 126 5502 900 5508
rect 1548 5508 1554 5511
rect 1548 5502 1584 5508
rect 126 5468 138 5502
rect 1572 5468 1584 5502
rect 126 5462 900 5468
rect 894 5459 900 5462
rect 1548 5462 1584 5468
rect 1548 5459 1554 5462
rect 156 5422 162 5425
rect 126 5416 162 5422
rect 810 5422 816 5425
rect 810 5416 1584 5422
rect 126 5382 138 5416
rect 1572 5382 1584 5416
rect 126 5376 162 5382
rect 156 5373 162 5376
rect 810 5376 1584 5382
rect 810 5373 816 5376
rect 894 5336 900 5339
rect 126 5330 900 5336
rect 1548 5336 1554 5339
rect 1548 5330 1584 5336
rect 126 5296 138 5330
rect 1572 5296 1584 5330
rect 126 5290 900 5296
rect 894 5287 900 5290
rect 1548 5290 1584 5296
rect 1548 5287 1554 5290
rect 156 5250 162 5253
rect 126 5244 162 5250
rect 810 5250 816 5253
rect 810 5244 1584 5250
rect 126 5210 138 5244
rect 1572 5210 1584 5244
rect 126 5204 162 5210
rect 156 5201 162 5204
rect 810 5204 1584 5210
rect 810 5201 816 5204
rect 894 5164 900 5167
rect 126 5158 900 5164
rect 1548 5164 1554 5167
rect 1548 5158 1584 5164
rect 126 5124 138 5158
rect 1572 5124 1584 5158
rect 126 5118 900 5124
rect 894 5115 900 5118
rect 1548 5118 1584 5124
rect 1548 5115 1554 5118
rect 156 5078 162 5081
rect 126 5072 162 5078
rect 810 5078 816 5081
rect 810 5072 1584 5078
rect 126 5038 138 5072
rect 1572 5038 1584 5072
rect 126 5032 162 5038
rect 156 5029 162 5032
rect 810 5032 1584 5038
rect 810 5029 816 5032
rect 894 4992 900 4995
rect 126 4986 900 4992
rect 1548 4992 1554 4995
rect 1548 4986 1584 4992
rect 126 4952 138 4986
rect 1572 4952 1584 4986
rect 126 4946 900 4952
rect 894 4943 900 4946
rect 1548 4946 1584 4952
rect 1548 4943 1554 4946
rect 156 4906 162 4909
rect 126 4900 162 4906
rect 810 4906 816 4909
rect 810 4900 1584 4906
rect 126 4866 138 4900
rect 1572 4866 1584 4900
rect 126 4860 162 4866
rect 156 4857 162 4860
rect 810 4860 1584 4866
rect 810 4857 816 4860
rect 894 4820 900 4823
rect 126 4814 900 4820
rect 1548 4820 1554 4823
rect 1548 4814 1584 4820
rect 126 4780 138 4814
rect 1572 4780 1584 4814
rect 126 4774 900 4780
rect 894 4771 900 4774
rect 1548 4774 1584 4780
rect 1548 4771 1554 4774
rect 156 4734 162 4737
rect 126 4728 162 4734
rect 810 4734 816 4737
rect 810 4728 1584 4734
rect 126 4694 138 4728
rect 1572 4694 1584 4728
rect 126 4688 162 4694
rect 156 4685 162 4688
rect 810 4688 1584 4694
rect 810 4685 816 4688
rect 894 4648 900 4651
rect 126 4642 900 4648
rect 1548 4648 1554 4651
rect 1548 4642 1584 4648
rect 126 4608 138 4642
rect 1572 4608 1584 4642
rect 126 4602 900 4608
rect 894 4599 900 4602
rect 1548 4602 1584 4608
rect 1548 4599 1554 4602
rect 156 4562 162 4565
rect 126 4556 162 4562
rect 810 4562 816 4565
rect 810 4556 1584 4562
rect 126 4522 138 4556
rect 1572 4522 1584 4556
rect 126 4516 162 4522
rect 156 4513 162 4516
rect 810 4516 1584 4522
rect 810 4513 816 4516
rect 894 4476 900 4479
rect 126 4470 900 4476
rect 1548 4476 1554 4479
rect 1548 4470 1584 4476
rect 126 4436 138 4470
rect 1572 4436 1584 4470
rect 126 4430 900 4436
rect 894 4427 900 4430
rect 1548 4430 1584 4436
rect 1548 4427 1554 4430
rect 156 4390 162 4393
rect 126 4384 162 4390
rect 810 4390 816 4393
rect 810 4384 1584 4390
rect 126 4350 138 4384
rect 1572 4350 1584 4384
rect 126 4344 162 4350
rect 156 4341 162 4344
rect 810 4344 1584 4350
rect 810 4341 816 4344
rect 894 4304 900 4307
rect 126 4298 900 4304
rect 1548 4304 1554 4307
rect 1548 4298 1584 4304
rect 126 4264 138 4298
rect 1572 4264 1584 4298
rect 126 4258 900 4264
rect 894 4255 900 4258
rect 1548 4258 1584 4264
rect 1548 4255 1554 4258
rect 156 4218 162 4221
rect 126 4212 162 4218
rect 810 4218 816 4221
rect 810 4212 1584 4218
rect 126 4178 138 4212
rect 1572 4178 1584 4212
rect 126 4172 162 4178
rect 156 4169 162 4172
rect 810 4172 1584 4178
rect 810 4169 816 4172
rect 894 4132 900 4135
rect 126 4126 900 4132
rect 1548 4132 1554 4135
rect 1548 4126 1584 4132
rect 126 4092 138 4126
rect 1572 4092 1584 4126
rect 126 4086 900 4092
rect 894 4083 900 4086
rect 1548 4086 1584 4092
rect 1548 4083 1554 4086
rect 156 4046 162 4049
rect 126 4040 162 4046
rect 810 4046 816 4049
rect 810 4040 1584 4046
rect 126 4006 138 4040
rect 1572 4006 1584 4040
rect 126 4000 162 4006
rect 156 3997 162 4000
rect 810 4000 1584 4006
rect 810 3997 816 4000
rect 894 3960 900 3963
rect 126 3954 900 3960
rect 1548 3960 1554 3963
rect 1548 3954 1584 3960
rect 126 3920 138 3954
rect 1572 3920 1584 3954
rect 126 3914 900 3920
rect 894 3911 900 3914
rect 1548 3914 1584 3920
rect 1548 3911 1554 3914
rect 156 3874 162 3877
rect 126 3868 162 3874
rect 810 3874 816 3877
rect 810 3868 1584 3874
rect 126 3834 138 3868
rect 1572 3834 1584 3868
rect 126 3828 162 3834
rect 156 3825 162 3828
rect 810 3828 1584 3834
rect 810 3825 816 3828
rect 894 3788 900 3791
rect 126 3782 900 3788
rect 1548 3788 1554 3791
rect 1548 3782 1584 3788
rect 126 3748 138 3782
rect 1572 3748 1584 3782
rect 126 3742 900 3748
rect 894 3739 900 3742
rect 1548 3742 1584 3748
rect 1548 3739 1554 3742
rect 156 3702 162 3705
rect 126 3696 162 3702
rect 810 3702 816 3705
rect 810 3696 1584 3702
rect 126 3662 138 3696
rect 1572 3662 1584 3696
rect 126 3656 162 3662
rect 156 3653 162 3656
rect 810 3656 1584 3662
rect 810 3653 816 3656
rect 894 3616 900 3619
rect 126 3610 900 3616
rect 1548 3616 1554 3619
rect 1548 3610 1584 3616
rect 126 3576 138 3610
rect 1572 3576 1584 3610
rect 126 3570 900 3576
rect 894 3567 900 3570
rect 1548 3570 1584 3576
rect 1548 3567 1554 3570
rect 156 3530 162 3533
rect 126 3524 162 3530
rect 810 3530 816 3533
rect 810 3524 1584 3530
rect 126 3490 138 3524
rect 1572 3490 1584 3524
rect 126 3484 162 3490
rect 156 3481 162 3484
rect 810 3484 1584 3490
rect 810 3481 816 3484
rect 894 3444 900 3447
rect 126 3438 900 3444
rect 1548 3444 1554 3447
rect 1548 3438 1584 3444
rect 126 3404 138 3438
rect 1572 3404 1584 3438
rect 126 3398 900 3404
rect 894 3395 900 3398
rect 1548 3398 1584 3404
rect 1548 3395 1554 3398
rect 156 3358 162 3361
rect 126 3352 162 3358
rect 810 3358 816 3361
rect 810 3352 1584 3358
rect 126 3318 138 3352
rect 1572 3318 1584 3352
rect 126 3312 162 3318
rect 156 3309 162 3312
rect 810 3312 1584 3318
rect 810 3309 816 3312
rect 894 3272 900 3275
rect 126 3266 900 3272
rect 1548 3272 1554 3275
rect 1548 3266 1584 3272
rect 126 3232 138 3266
rect 1572 3232 1584 3266
rect 126 3226 900 3232
rect 894 3223 900 3226
rect 1548 3226 1584 3232
rect 1548 3223 1554 3226
rect 156 3186 162 3189
rect 126 3180 162 3186
rect 810 3186 816 3189
rect 810 3180 1584 3186
rect 126 3146 138 3180
rect 1572 3146 1584 3180
rect 126 3140 162 3146
rect 156 3137 162 3140
rect 810 3140 1584 3146
rect 810 3137 816 3140
rect 894 3100 900 3103
rect 126 3094 900 3100
rect 1548 3100 1554 3103
rect 1548 3094 1584 3100
rect 126 3060 138 3094
rect 1572 3060 1584 3094
rect 126 3054 900 3060
rect 894 3051 900 3054
rect 1548 3054 1584 3060
rect 1548 3051 1554 3054
rect 156 3014 162 3017
rect 126 3008 162 3014
rect 810 3014 816 3017
rect 810 3008 1584 3014
rect 126 2974 138 3008
rect 1572 2974 1584 3008
rect 126 2968 162 2974
rect 156 2965 162 2968
rect 810 2968 1584 2974
rect 810 2965 816 2968
rect 894 2928 900 2931
rect 126 2922 900 2928
rect 1548 2928 1554 2931
rect 1548 2922 1584 2928
rect 126 2888 138 2922
rect 1572 2888 1584 2922
rect 126 2882 900 2888
rect 894 2879 900 2882
rect 1548 2882 1584 2888
rect 1548 2879 1554 2882
rect 156 2842 162 2845
rect 126 2836 162 2842
rect 810 2842 816 2845
rect 810 2836 1584 2842
rect 126 2802 138 2836
rect 1572 2802 1584 2836
rect 126 2796 162 2802
rect 156 2793 162 2796
rect 810 2796 1584 2802
rect 810 2793 816 2796
rect 894 2756 900 2759
rect 126 2750 900 2756
rect 1548 2756 1554 2759
rect 1548 2750 1584 2756
rect 126 2716 138 2750
rect 1572 2716 1584 2750
rect 126 2710 900 2716
rect 894 2707 900 2710
rect 1548 2710 1584 2716
rect 1548 2707 1554 2710
rect 156 2670 162 2673
rect 126 2664 162 2670
rect 810 2670 816 2673
rect 810 2664 1584 2670
rect 126 2630 138 2664
rect 1572 2630 1584 2664
rect 126 2624 162 2630
rect 156 2621 162 2624
rect 810 2624 1584 2630
rect 810 2621 816 2624
rect 894 2584 900 2587
rect 126 2578 900 2584
rect 1548 2584 1554 2587
rect 1548 2578 1584 2584
rect 126 2544 138 2578
rect 1572 2544 1584 2578
rect 126 2538 900 2544
rect 894 2535 900 2538
rect 1548 2538 1584 2544
rect 1548 2535 1554 2538
rect 156 2498 162 2501
rect 126 2492 162 2498
rect 810 2498 816 2501
rect 810 2492 1584 2498
rect 126 2458 138 2492
rect 1572 2458 1584 2492
rect 126 2452 162 2458
rect 156 2449 162 2452
rect 810 2452 1584 2458
rect 810 2449 816 2452
rect 894 2412 900 2415
rect 126 2406 900 2412
rect 1548 2412 1554 2415
rect 1548 2406 1584 2412
rect 126 2372 138 2406
rect 1572 2372 1584 2406
rect 126 2366 900 2372
rect 894 2363 900 2366
rect 1548 2366 1584 2372
rect 1548 2363 1554 2366
rect 156 2326 162 2329
rect 126 2320 162 2326
rect 810 2326 816 2329
rect 810 2320 1584 2326
rect 126 2286 138 2320
rect 1572 2286 1584 2320
rect 126 2280 162 2286
rect 156 2277 162 2280
rect 810 2280 1584 2286
rect 810 2277 816 2280
rect 894 2240 900 2243
rect 126 2234 900 2240
rect 1548 2240 1554 2243
rect 1548 2234 1584 2240
rect 126 2200 138 2234
rect 1572 2200 1584 2234
rect 126 2194 900 2200
rect 894 2191 900 2194
rect 1548 2194 1584 2200
rect 1548 2191 1554 2194
rect 156 2154 162 2157
rect 126 2148 162 2154
rect 810 2154 816 2157
rect 810 2148 1584 2154
rect 126 2114 138 2148
rect 1572 2114 1584 2148
rect 126 2108 162 2114
rect 156 2105 162 2108
rect 810 2108 1584 2114
rect 810 2105 816 2108
rect 894 2068 900 2071
rect 126 2062 900 2068
rect 1548 2068 1554 2071
rect 1548 2062 1584 2068
rect 126 2028 138 2062
rect 1572 2028 1584 2062
rect 126 2022 900 2028
rect 894 2019 900 2022
rect 1548 2022 1584 2028
rect 1548 2019 1554 2022
rect 156 1982 162 1985
rect 126 1976 162 1982
rect 810 1982 816 1985
rect 810 1976 1584 1982
rect 126 1942 138 1976
rect 1572 1942 1584 1976
rect 126 1936 162 1942
rect 156 1933 162 1936
rect 810 1936 1584 1942
rect 810 1933 816 1936
rect 894 1896 900 1899
rect 126 1890 900 1896
rect 1548 1896 1554 1899
rect 1548 1890 1584 1896
rect 126 1856 138 1890
rect 1572 1856 1584 1890
rect 126 1850 900 1856
rect 894 1847 900 1850
rect 1548 1850 1584 1856
rect 1548 1847 1554 1850
rect 156 1810 162 1813
rect 126 1804 162 1810
rect 810 1810 816 1813
rect 810 1804 1584 1810
rect 126 1770 138 1804
rect 1572 1770 1584 1804
rect 126 1764 162 1770
rect 156 1761 162 1764
rect 810 1764 1584 1770
rect 810 1761 816 1764
rect 894 1724 900 1727
rect 126 1718 900 1724
rect 1548 1724 1554 1727
rect 1548 1718 1584 1724
rect 126 1684 138 1718
rect 1572 1684 1584 1718
rect 126 1678 900 1684
rect 894 1675 900 1678
rect 1548 1678 1584 1684
rect 1548 1675 1554 1678
rect 156 1638 162 1641
rect 126 1632 162 1638
rect 810 1638 816 1641
rect 810 1632 1584 1638
rect 126 1598 138 1632
rect 1572 1598 1584 1632
rect 126 1592 162 1598
rect 156 1589 162 1592
rect 810 1592 1584 1598
rect 810 1589 816 1592
rect 894 1552 900 1555
rect 126 1546 900 1552
rect 1548 1552 1554 1555
rect 1548 1546 1584 1552
rect 126 1512 138 1546
rect 1572 1512 1584 1546
rect 126 1506 900 1512
rect 894 1503 900 1506
rect 1548 1506 1584 1512
rect 1548 1503 1554 1506
rect 156 1466 162 1469
rect 126 1460 162 1466
rect 810 1466 816 1469
rect 810 1460 1584 1466
rect 126 1426 138 1460
rect 1572 1426 1584 1460
rect 126 1420 162 1426
rect 156 1417 162 1420
rect 810 1420 1584 1426
rect 810 1417 816 1420
rect 894 1380 900 1383
rect 126 1374 900 1380
rect 1548 1380 1554 1383
rect 1548 1374 1584 1380
rect 126 1340 138 1374
rect 1572 1340 1584 1374
rect 126 1334 900 1340
rect 894 1331 900 1334
rect 1548 1334 1584 1340
rect 1548 1331 1554 1334
rect 156 1294 162 1297
rect 126 1288 162 1294
rect 810 1294 816 1297
rect 810 1288 1584 1294
rect 126 1254 138 1288
rect 1572 1254 1584 1288
rect 126 1248 162 1254
rect 156 1245 162 1248
rect 810 1248 1584 1254
rect 810 1245 816 1248
rect 894 1208 900 1211
rect 126 1202 900 1208
rect 1548 1208 1554 1211
rect 1548 1202 1584 1208
rect 126 1168 138 1202
rect 1572 1168 1584 1202
rect 126 1162 900 1168
rect 894 1159 900 1162
rect 1548 1162 1584 1168
rect 1548 1159 1554 1162
rect 156 1122 162 1125
rect 126 1116 162 1122
rect 810 1122 816 1125
rect 810 1116 1584 1122
rect 126 1082 138 1116
rect 1572 1082 1584 1116
rect 126 1076 162 1082
rect 156 1073 162 1076
rect 810 1076 1584 1082
rect 810 1073 816 1076
rect 894 1036 900 1039
rect 126 1030 900 1036
rect 1548 1036 1554 1039
rect 1548 1030 1584 1036
rect 126 996 138 1030
rect 1572 996 1584 1030
rect 126 990 900 996
rect 894 987 900 990
rect 1548 990 1584 996
rect 1548 987 1554 990
rect 156 950 162 953
rect 126 944 162 950
rect 810 950 816 953
rect 810 944 1584 950
rect 126 910 138 944
rect 1572 910 1584 944
rect 126 904 162 910
rect 156 901 162 904
rect 810 904 1584 910
rect 810 901 816 904
rect 894 864 900 867
rect 126 858 900 864
rect 1548 864 1554 867
rect 1548 858 1584 864
rect 126 824 138 858
rect 1572 824 1584 858
rect 126 818 900 824
rect 894 815 900 818
rect 1548 818 1584 824
rect 1548 815 1554 818
rect 156 778 162 781
rect 126 772 162 778
rect 810 778 816 781
rect 810 772 1584 778
rect 126 738 138 772
rect 1572 738 1584 772
rect 126 732 162 738
rect 156 729 162 732
rect 810 732 1584 738
rect 810 729 816 732
rect 894 692 900 695
rect 126 686 900 692
rect 1548 692 1554 695
rect 1548 686 1584 692
rect 126 652 138 686
rect 1572 652 1584 686
rect 126 646 900 652
rect 894 643 900 646
rect 1548 646 1584 652
rect 1548 643 1554 646
rect 156 606 162 609
rect 126 600 162 606
rect 810 606 816 609
rect 810 600 1584 606
rect 126 566 138 600
rect 1572 566 1584 600
rect 126 560 162 566
rect 156 557 162 560
rect 810 560 1584 566
rect 810 557 816 560
rect 894 520 900 523
rect 126 514 900 520
rect 1548 520 1554 523
rect 1548 514 1584 520
rect 126 480 138 514
rect 1572 480 1584 514
rect 126 474 900 480
rect 894 471 900 474
rect 1548 474 1584 480
rect 1548 471 1554 474
rect 156 434 162 437
rect 126 428 162 434
rect 810 434 816 437
rect 810 428 1584 434
rect 126 394 138 428
rect 1572 394 1584 428
rect 126 388 162 394
rect 156 385 162 388
rect 810 388 1584 394
rect 810 385 816 388
rect 894 348 900 351
rect 126 342 900 348
rect 1548 348 1554 351
rect 1548 342 1584 348
rect 126 308 138 342
rect 1572 308 1584 342
rect 126 302 900 308
rect 894 299 900 302
rect 1548 302 1584 308
rect 1548 299 1554 302
rect 156 262 162 265
rect 126 256 162 262
rect 810 262 816 265
rect 810 256 1584 262
rect 126 222 138 256
rect 1572 222 1584 256
rect 126 216 162 222
rect 156 213 162 216
rect 810 216 1584 222
rect 810 213 816 216
rect 894 176 900 179
rect 126 170 900 176
rect 1548 176 1554 179
rect 1548 170 1584 176
rect 126 136 138 170
rect 1572 136 1584 170
rect 1618 163 1672 169
rect 126 130 900 136
rect 894 127 900 130
rect 1548 130 1584 136
rect 1548 127 1554 130
rect 30 76 76 100
rect 1704 100 1710 43894
rect 1744 100 1750 43894
rect 1704 76 1750 100
rect 30 70 1750 76
rect 30 36 100 70
rect 1680 36 1750 70
rect 30 30 1750 36
<< via1 >>
rect 900 43858 1548 43867
rect 900 43824 1548 43858
rect 900 43815 1548 43824
rect 1618 43815 1672 43825
rect 162 43772 810 43781
rect 162 43738 810 43772
rect 162 43729 810 43738
rect 900 43686 1548 43695
rect 900 43652 1548 43686
rect 900 43643 1548 43652
rect 162 43600 810 43609
rect 162 43566 810 43600
rect 162 43557 810 43566
rect 900 43514 1548 43523
rect 900 43480 1548 43514
rect 900 43471 1548 43480
rect 162 43428 810 43437
rect 162 43394 810 43428
rect 162 43385 810 43394
rect 900 43342 1548 43351
rect 900 43308 1548 43342
rect 900 43299 1548 43308
rect 162 43256 810 43265
rect 162 43222 810 43256
rect 162 43213 810 43222
rect 900 43170 1548 43179
rect 900 43136 1548 43170
rect 900 43127 1548 43136
rect 162 43084 810 43093
rect 162 43050 810 43084
rect 162 43041 810 43050
rect 900 42998 1548 43007
rect 900 42964 1548 42998
rect 900 42955 1548 42964
rect 162 42912 810 42921
rect 162 42878 810 42912
rect 162 42869 810 42878
rect 900 42826 1548 42835
rect 900 42792 1548 42826
rect 900 42783 1548 42792
rect 162 42740 810 42749
rect 162 42706 810 42740
rect 162 42697 810 42706
rect 900 42654 1548 42663
rect 900 42620 1548 42654
rect 900 42611 1548 42620
rect 162 42568 810 42577
rect 162 42534 810 42568
rect 162 42525 810 42534
rect 900 42482 1548 42491
rect 900 42448 1548 42482
rect 900 42439 1548 42448
rect 162 42396 810 42405
rect 162 42362 810 42396
rect 162 42353 810 42362
rect 900 42310 1548 42319
rect 900 42276 1548 42310
rect 900 42267 1548 42276
rect 162 42224 810 42233
rect 162 42190 810 42224
rect 162 42181 810 42190
rect 900 42138 1548 42147
rect 900 42104 1548 42138
rect 900 42095 1548 42104
rect 162 42052 810 42061
rect 162 42018 810 42052
rect 162 42009 810 42018
rect 900 41966 1548 41975
rect 900 41932 1548 41966
rect 900 41923 1548 41932
rect 162 41880 810 41889
rect 162 41846 810 41880
rect 162 41837 810 41846
rect 900 41794 1548 41803
rect 900 41760 1548 41794
rect 900 41751 1548 41760
rect 162 41708 810 41717
rect 162 41674 810 41708
rect 162 41665 810 41674
rect 900 41622 1548 41631
rect 900 41588 1548 41622
rect 900 41579 1548 41588
rect 162 41536 810 41545
rect 162 41502 810 41536
rect 162 41493 810 41502
rect 900 41450 1548 41459
rect 900 41416 1548 41450
rect 900 41407 1548 41416
rect 162 41364 810 41373
rect 162 41330 810 41364
rect 162 41321 810 41330
rect 900 41278 1548 41287
rect 900 41244 1548 41278
rect 900 41235 1548 41244
rect 162 41192 810 41201
rect 162 41158 810 41192
rect 162 41149 810 41158
rect 900 41106 1548 41115
rect 900 41072 1548 41106
rect 900 41063 1548 41072
rect 162 41020 810 41029
rect 162 40986 810 41020
rect 162 40977 810 40986
rect 900 40934 1548 40943
rect 900 40900 1548 40934
rect 900 40891 1548 40900
rect 162 40848 810 40857
rect 162 40814 810 40848
rect 162 40805 810 40814
rect 900 40762 1548 40771
rect 900 40728 1548 40762
rect 900 40719 1548 40728
rect 162 40676 810 40685
rect 162 40642 810 40676
rect 162 40633 810 40642
rect 900 40590 1548 40599
rect 900 40556 1548 40590
rect 900 40547 1548 40556
rect 162 40504 810 40513
rect 162 40470 810 40504
rect 162 40461 810 40470
rect 900 40418 1548 40427
rect 900 40384 1548 40418
rect 900 40375 1548 40384
rect 162 40332 810 40341
rect 162 40298 810 40332
rect 162 40289 810 40298
rect 900 40246 1548 40255
rect 900 40212 1548 40246
rect 900 40203 1548 40212
rect 162 40160 810 40169
rect 162 40126 810 40160
rect 162 40117 810 40126
rect 900 40074 1548 40083
rect 900 40040 1548 40074
rect 900 40031 1548 40040
rect 162 39988 810 39997
rect 162 39954 810 39988
rect 162 39945 810 39954
rect 900 39902 1548 39911
rect 900 39868 1548 39902
rect 900 39859 1548 39868
rect 162 39816 810 39825
rect 162 39782 810 39816
rect 162 39773 810 39782
rect 900 39730 1548 39739
rect 900 39696 1548 39730
rect 900 39687 1548 39696
rect 162 39644 810 39653
rect 162 39610 810 39644
rect 162 39601 810 39610
rect 900 39558 1548 39567
rect 900 39524 1548 39558
rect 900 39515 1548 39524
rect 162 39472 810 39481
rect 162 39438 810 39472
rect 162 39429 810 39438
rect 900 39386 1548 39395
rect 900 39352 1548 39386
rect 900 39343 1548 39352
rect 162 39300 810 39309
rect 162 39266 810 39300
rect 162 39257 810 39266
rect 900 39214 1548 39223
rect 900 39180 1548 39214
rect 900 39171 1548 39180
rect 162 39128 810 39137
rect 162 39094 810 39128
rect 162 39085 810 39094
rect 900 39042 1548 39051
rect 900 39008 1548 39042
rect 900 38999 1548 39008
rect 162 38956 810 38965
rect 162 38922 810 38956
rect 162 38913 810 38922
rect 900 38870 1548 38879
rect 900 38836 1548 38870
rect 900 38827 1548 38836
rect 162 38784 810 38793
rect 162 38750 810 38784
rect 162 38741 810 38750
rect 900 38698 1548 38707
rect 900 38664 1548 38698
rect 900 38655 1548 38664
rect 162 38612 810 38621
rect 162 38578 810 38612
rect 162 38569 810 38578
rect 900 38526 1548 38535
rect 900 38492 1548 38526
rect 900 38483 1548 38492
rect 162 38440 810 38449
rect 162 38406 810 38440
rect 162 38397 810 38406
rect 900 38354 1548 38363
rect 900 38320 1548 38354
rect 900 38311 1548 38320
rect 162 38268 810 38277
rect 162 38234 810 38268
rect 162 38225 810 38234
rect 900 38182 1548 38191
rect 900 38148 1548 38182
rect 900 38139 1548 38148
rect 162 38096 810 38105
rect 162 38062 810 38096
rect 162 38053 810 38062
rect 900 38010 1548 38019
rect 900 37976 1548 38010
rect 900 37967 1548 37976
rect 162 37924 810 37933
rect 162 37890 810 37924
rect 162 37881 810 37890
rect 900 37838 1548 37847
rect 900 37804 1548 37838
rect 900 37795 1548 37804
rect 162 37752 810 37761
rect 162 37718 810 37752
rect 162 37709 810 37718
rect 900 37666 1548 37675
rect 900 37632 1548 37666
rect 900 37623 1548 37632
rect 162 37580 810 37589
rect 162 37546 810 37580
rect 162 37537 810 37546
rect 900 37494 1548 37503
rect 900 37460 1548 37494
rect 900 37451 1548 37460
rect 162 37408 810 37417
rect 162 37374 810 37408
rect 162 37365 810 37374
rect 900 37322 1548 37331
rect 900 37288 1548 37322
rect 900 37279 1548 37288
rect 162 37236 810 37245
rect 162 37202 810 37236
rect 162 37193 810 37202
rect 900 37150 1548 37159
rect 900 37116 1548 37150
rect 900 37107 1548 37116
rect 162 37064 810 37073
rect 162 37030 810 37064
rect 162 37021 810 37030
rect 900 36978 1548 36987
rect 900 36944 1548 36978
rect 900 36935 1548 36944
rect 162 36892 810 36901
rect 162 36858 810 36892
rect 162 36849 810 36858
rect 900 36806 1548 36815
rect 900 36772 1548 36806
rect 900 36763 1548 36772
rect 162 36720 810 36729
rect 162 36686 810 36720
rect 162 36677 810 36686
rect 900 36634 1548 36643
rect 900 36600 1548 36634
rect 900 36591 1548 36600
rect 162 36548 810 36557
rect 162 36514 810 36548
rect 162 36505 810 36514
rect 900 36462 1548 36471
rect 900 36428 1548 36462
rect 900 36419 1548 36428
rect 162 36376 810 36385
rect 162 36342 810 36376
rect 162 36333 810 36342
rect 900 36290 1548 36299
rect 900 36256 1548 36290
rect 900 36247 1548 36256
rect 162 36204 810 36213
rect 162 36170 810 36204
rect 162 36161 810 36170
rect 900 36118 1548 36127
rect 900 36084 1548 36118
rect 900 36075 1548 36084
rect 162 36032 810 36041
rect 162 35998 810 36032
rect 162 35989 810 35998
rect 900 35946 1548 35955
rect 900 35912 1548 35946
rect 900 35903 1548 35912
rect 162 35860 810 35869
rect 162 35826 810 35860
rect 162 35817 810 35826
rect 900 35774 1548 35783
rect 900 35740 1548 35774
rect 900 35731 1548 35740
rect 162 35688 810 35697
rect 162 35654 810 35688
rect 162 35645 810 35654
rect 900 35602 1548 35611
rect 900 35568 1548 35602
rect 900 35559 1548 35568
rect 162 35516 810 35525
rect 162 35482 810 35516
rect 162 35473 810 35482
rect 900 35430 1548 35439
rect 900 35396 1548 35430
rect 900 35387 1548 35396
rect 162 35344 810 35353
rect 162 35310 810 35344
rect 162 35301 810 35310
rect 900 35258 1548 35267
rect 900 35224 1548 35258
rect 900 35215 1548 35224
rect 162 35172 810 35181
rect 162 35138 810 35172
rect 162 35129 810 35138
rect 900 35086 1548 35095
rect 900 35052 1548 35086
rect 900 35043 1548 35052
rect 162 35000 810 35009
rect 162 34966 810 35000
rect 162 34957 810 34966
rect 900 34914 1548 34923
rect 900 34880 1548 34914
rect 900 34871 1548 34880
rect 162 34828 810 34837
rect 162 34794 810 34828
rect 162 34785 810 34794
rect 900 34742 1548 34751
rect 900 34708 1548 34742
rect 900 34699 1548 34708
rect 162 34656 810 34665
rect 162 34622 810 34656
rect 162 34613 810 34622
rect 900 34570 1548 34579
rect 900 34536 1548 34570
rect 900 34527 1548 34536
rect 162 34484 810 34493
rect 162 34450 810 34484
rect 162 34441 810 34450
rect 900 34398 1548 34407
rect 900 34364 1548 34398
rect 900 34355 1548 34364
rect 162 34312 810 34321
rect 162 34278 810 34312
rect 162 34269 810 34278
rect 900 34226 1548 34235
rect 900 34192 1548 34226
rect 900 34183 1548 34192
rect 162 34140 810 34149
rect 162 34106 810 34140
rect 162 34097 810 34106
rect 900 34054 1548 34063
rect 900 34020 1548 34054
rect 900 34011 1548 34020
rect 162 33968 810 33977
rect 162 33934 810 33968
rect 162 33925 810 33934
rect 900 33882 1548 33891
rect 900 33848 1548 33882
rect 900 33839 1548 33848
rect 162 33796 810 33805
rect 162 33762 810 33796
rect 162 33753 810 33762
rect 900 33710 1548 33719
rect 900 33676 1548 33710
rect 900 33667 1548 33676
rect 162 33624 810 33633
rect 162 33590 810 33624
rect 162 33581 810 33590
rect 900 33538 1548 33547
rect 900 33504 1548 33538
rect 900 33495 1548 33504
rect 162 33452 810 33461
rect 162 33418 810 33452
rect 162 33409 810 33418
rect 900 33366 1548 33375
rect 900 33332 1548 33366
rect 900 33323 1548 33332
rect 162 33280 810 33289
rect 162 33246 810 33280
rect 162 33237 810 33246
rect 900 33194 1548 33203
rect 900 33160 1548 33194
rect 900 33151 1548 33160
rect 162 33108 810 33117
rect 162 33074 810 33108
rect 162 33065 810 33074
rect 900 33022 1548 33031
rect 900 32988 1548 33022
rect 900 32979 1548 32988
rect 162 32936 810 32945
rect 162 32902 810 32936
rect 162 32893 810 32902
rect 900 32850 1548 32859
rect 900 32816 1548 32850
rect 900 32807 1548 32816
rect 162 32764 810 32773
rect 162 32730 810 32764
rect 162 32721 810 32730
rect 900 32678 1548 32687
rect 900 32644 1548 32678
rect 900 32635 1548 32644
rect 162 32592 810 32601
rect 162 32558 810 32592
rect 162 32549 810 32558
rect 900 32506 1548 32515
rect 900 32472 1548 32506
rect 900 32463 1548 32472
rect 162 32420 810 32429
rect 162 32386 810 32420
rect 162 32377 810 32386
rect 900 32334 1548 32343
rect 900 32300 1548 32334
rect 900 32291 1548 32300
rect 162 32248 810 32257
rect 162 32214 810 32248
rect 162 32205 810 32214
rect 900 32162 1548 32171
rect 900 32128 1548 32162
rect 900 32119 1548 32128
rect 162 32076 810 32085
rect 162 32042 810 32076
rect 162 32033 810 32042
rect 900 31990 1548 31999
rect 900 31956 1548 31990
rect 900 31947 1548 31956
rect 162 31904 810 31913
rect 162 31870 810 31904
rect 162 31861 810 31870
rect 900 31818 1548 31827
rect 900 31784 1548 31818
rect 900 31775 1548 31784
rect 162 31732 810 31741
rect 162 31698 810 31732
rect 162 31689 810 31698
rect 900 31646 1548 31655
rect 900 31612 1548 31646
rect 900 31603 1548 31612
rect 162 31560 810 31569
rect 162 31526 810 31560
rect 162 31517 810 31526
rect 900 31474 1548 31483
rect 900 31440 1548 31474
rect 900 31431 1548 31440
rect 162 31388 810 31397
rect 162 31354 810 31388
rect 162 31345 810 31354
rect 900 31302 1548 31311
rect 900 31268 1548 31302
rect 900 31259 1548 31268
rect 162 31216 810 31225
rect 162 31182 810 31216
rect 162 31173 810 31182
rect 900 31130 1548 31139
rect 900 31096 1548 31130
rect 900 31087 1548 31096
rect 162 31044 810 31053
rect 162 31010 810 31044
rect 162 31001 810 31010
rect 900 30958 1548 30967
rect 900 30924 1548 30958
rect 900 30915 1548 30924
rect 162 30872 810 30881
rect 162 30838 810 30872
rect 162 30829 810 30838
rect 900 30786 1548 30795
rect 900 30752 1548 30786
rect 900 30743 1548 30752
rect 162 30700 810 30709
rect 162 30666 810 30700
rect 162 30657 810 30666
rect 900 30614 1548 30623
rect 900 30580 1548 30614
rect 900 30571 1548 30580
rect 162 30528 810 30537
rect 162 30494 810 30528
rect 162 30485 810 30494
rect 900 30442 1548 30451
rect 900 30408 1548 30442
rect 900 30399 1548 30408
rect 162 30356 810 30365
rect 162 30322 810 30356
rect 162 30313 810 30322
rect 900 30270 1548 30279
rect 900 30236 1548 30270
rect 900 30227 1548 30236
rect 162 30184 810 30193
rect 162 30150 810 30184
rect 162 30141 810 30150
rect 900 30098 1548 30107
rect 900 30064 1548 30098
rect 900 30055 1548 30064
rect 162 30012 810 30021
rect 162 29978 810 30012
rect 162 29969 810 29978
rect 900 29926 1548 29935
rect 900 29892 1548 29926
rect 900 29883 1548 29892
rect 162 29840 810 29849
rect 162 29806 810 29840
rect 162 29797 810 29806
rect 900 29754 1548 29763
rect 900 29720 1548 29754
rect 900 29711 1548 29720
rect 162 29668 810 29677
rect 162 29634 810 29668
rect 162 29625 810 29634
rect 900 29582 1548 29591
rect 900 29548 1548 29582
rect 900 29539 1548 29548
rect 162 29496 810 29505
rect 162 29462 810 29496
rect 162 29453 810 29462
rect 900 29410 1548 29419
rect 900 29376 1548 29410
rect 900 29367 1548 29376
rect 162 29324 810 29333
rect 162 29290 810 29324
rect 162 29281 810 29290
rect 900 29238 1548 29247
rect 900 29204 1548 29238
rect 900 29195 1548 29204
rect 162 29152 810 29161
rect 162 29118 810 29152
rect 162 29109 810 29118
rect 900 29066 1548 29075
rect 900 29032 1548 29066
rect 900 29023 1548 29032
rect 162 28980 810 28989
rect 162 28946 810 28980
rect 162 28937 810 28946
rect 900 28894 1548 28903
rect 900 28860 1548 28894
rect 900 28851 1548 28860
rect 162 28808 810 28817
rect 162 28774 810 28808
rect 162 28765 810 28774
rect 900 28722 1548 28731
rect 900 28688 1548 28722
rect 900 28679 1548 28688
rect 162 28636 810 28645
rect 162 28602 810 28636
rect 162 28593 810 28602
rect 900 28550 1548 28559
rect 900 28516 1548 28550
rect 900 28507 1548 28516
rect 162 28464 810 28473
rect 162 28430 810 28464
rect 162 28421 810 28430
rect 900 28378 1548 28387
rect 900 28344 1548 28378
rect 900 28335 1548 28344
rect 162 28292 810 28301
rect 162 28258 810 28292
rect 162 28249 810 28258
rect 900 28206 1548 28215
rect 900 28172 1548 28206
rect 900 28163 1548 28172
rect 162 28120 810 28129
rect 162 28086 810 28120
rect 162 28077 810 28086
rect 900 28034 1548 28043
rect 900 28000 1548 28034
rect 900 27991 1548 28000
rect 162 27948 810 27957
rect 162 27914 810 27948
rect 162 27905 810 27914
rect 900 27862 1548 27871
rect 900 27828 1548 27862
rect 900 27819 1548 27828
rect 162 27776 810 27785
rect 162 27742 810 27776
rect 162 27733 810 27742
rect 900 27690 1548 27699
rect 900 27656 1548 27690
rect 900 27647 1548 27656
rect 162 27604 810 27613
rect 162 27570 810 27604
rect 162 27561 810 27570
rect 900 27518 1548 27527
rect 900 27484 1548 27518
rect 900 27475 1548 27484
rect 162 27432 810 27441
rect 162 27398 810 27432
rect 162 27389 810 27398
rect 900 27346 1548 27355
rect 900 27312 1548 27346
rect 900 27303 1548 27312
rect 162 27260 810 27269
rect 162 27226 810 27260
rect 162 27217 810 27226
rect 900 27174 1548 27183
rect 900 27140 1548 27174
rect 900 27131 1548 27140
rect 162 27088 810 27097
rect 162 27054 810 27088
rect 162 27045 810 27054
rect 900 27002 1548 27011
rect 900 26968 1548 27002
rect 900 26959 1548 26968
rect 162 26916 810 26925
rect 162 26882 810 26916
rect 162 26873 810 26882
rect 900 26830 1548 26839
rect 900 26796 1548 26830
rect 900 26787 1548 26796
rect 162 26744 810 26753
rect 162 26710 810 26744
rect 162 26701 810 26710
rect 900 26658 1548 26667
rect 900 26624 1548 26658
rect 900 26615 1548 26624
rect 162 26572 810 26581
rect 162 26538 810 26572
rect 162 26529 810 26538
rect 900 26486 1548 26495
rect 900 26452 1548 26486
rect 900 26443 1548 26452
rect 162 26400 810 26409
rect 162 26366 810 26400
rect 162 26357 810 26366
rect 900 26314 1548 26323
rect 900 26280 1548 26314
rect 900 26271 1548 26280
rect 162 26228 810 26237
rect 162 26194 810 26228
rect 162 26185 810 26194
rect 900 26142 1548 26151
rect 900 26108 1548 26142
rect 900 26099 1548 26108
rect 162 26056 810 26065
rect 162 26022 810 26056
rect 162 26013 810 26022
rect 900 25970 1548 25979
rect 900 25936 1548 25970
rect 900 25927 1548 25936
rect 162 25884 810 25893
rect 162 25850 810 25884
rect 162 25841 810 25850
rect 900 25798 1548 25807
rect 900 25764 1548 25798
rect 900 25755 1548 25764
rect 162 25712 810 25721
rect 162 25678 810 25712
rect 162 25669 810 25678
rect 900 25626 1548 25635
rect 900 25592 1548 25626
rect 900 25583 1548 25592
rect 162 25540 810 25549
rect 162 25506 810 25540
rect 162 25497 810 25506
rect 900 25454 1548 25463
rect 900 25420 1548 25454
rect 900 25411 1548 25420
rect 162 25368 810 25377
rect 162 25334 810 25368
rect 162 25325 810 25334
rect 900 25282 1548 25291
rect 900 25248 1548 25282
rect 900 25239 1548 25248
rect 162 25196 810 25205
rect 162 25162 810 25196
rect 162 25153 810 25162
rect 900 25110 1548 25119
rect 900 25076 1548 25110
rect 900 25067 1548 25076
rect 162 25024 810 25033
rect 162 24990 810 25024
rect 162 24981 810 24990
rect 900 24938 1548 24947
rect 900 24904 1548 24938
rect 900 24895 1548 24904
rect 162 24852 810 24861
rect 162 24818 810 24852
rect 162 24809 810 24818
rect 900 24766 1548 24775
rect 900 24732 1548 24766
rect 900 24723 1548 24732
rect 162 24680 810 24689
rect 162 24646 810 24680
rect 162 24637 810 24646
rect 900 24594 1548 24603
rect 900 24560 1548 24594
rect 900 24551 1548 24560
rect 162 24508 810 24517
rect 162 24474 810 24508
rect 162 24465 810 24474
rect 900 24422 1548 24431
rect 900 24388 1548 24422
rect 900 24379 1548 24388
rect 162 24336 810 24345
rect 162 24302 810 24336
rect 162 24293 810 24302
rect 900 24250 1548 24259
rect 900 24216 1548 24250
rect 900 24207 1548 24216
rect 162 24164 810 24173
rect 162 24130 810 24164
rect 162 24121 810 24130
rect 900 24078 1548 24087
rect 900 24044 1548 24078
rect 900 24035 1548 24044
rect 162 23992 810 24001
rect 162 23958 810 23992
rect 162 23949 810 23958
rect 900 23906 1548 23915
rect 900 23872 1548 23906
rect 900 23863 1548 23872
rect 162 23820 810 23829
rect 162 23786 810 23820
rect 162 23777 810 23786
rect 900 23734 1548 23743
rect 900 23700 1548 23734
rect 900 23691 1548 23700
rect 162 23648 810 23657
rect 162 23614 810 23648
rect 162 23605 810 23614
rect 900 23562 1548 23571
rect 900 23528 1548 23562
rect 900 23519 1548 23528
rect 162 23476 810 23485
rect 162 23442 810 23476
rect 162 23433 810 23442
rect 900 23390 1548 23399
rect 900 23356 1548 23390
rect 900 23347 1548 23356
rect 162 23304 810 23313
rect 162 23270 810 23304
rect 162 23261 810 23270
rect 900 23218 1548 23227
rect 900 23184 1548 23218
rect 900 23175 1548 23184
rect 162 23132 810 23141
rect 162 23098 810 23132
rect 162 23089 810 23098
rect 900 23046 1548 23055
rect 900 23012 1548 23046
rect 900 23003 1548 23012
rect 162 22960 810 22969
rect 162 22926 810 22960
rect 162 22917 810 22926
rect 900 22874 1548 22883
rect 900 22840 1548 22874
rect 900 22831 1548 22840
rect 162 22788 810 22797
rect 162 22754 810 22788
rect 162 22745 810 22754
rect 900 22702 1548 22711
rect 900 22668 1548 22702
rect 900 22659 1548 22668
rect 162 22616 810 22625
rect 162 22582 810 22616
rect 162 22573 810 22582
rect 900 22530 1548 22539
rect 900 22496 1548 22530
rect 900 22487 1548 22496
rect 162 22444 810 22453
rect 162 22410 810 22444
rect 162 22401 810 22410
rect 900 22358 1548 22367
rect 900 22324 1548 22358
rect 900 22315 1548 22324
rect 162 22272 810 22281
rect 162 22238 810 22272
rect 162 22229 810 22238
rect 900 22186 1548 22195
rect 900 22152 1548 22186
rect 900 22143 1548 22152
rect 162 22100 810 22109
rect 162 22066 810 22100
rect 162 22057 810 22066
rect 900 22014 1548 22023
rect 900 21980 1548 22014
rect 900 21971 1548 21980
rect 162 21928 810 21937
rect 162 21894 810 21928
rect 162 21885 810 21894
rect 900 21842 1548 21851
rect 900 21808 1548 21842
rect 900 21799 1548 21808
rect 162 21756 810 21765
rect 162 21722 810 21756
rect 162 21713 810 21722
rect 900 21670 1548 21679
rect 900 21636 1548 21670
rect 900 21627 1548 21636
rect 162 21584 810 21593
rect 162 21550 810 21584
rect 162 21541 810 21550
rect 900 21498 1548 21507
rect 900 21464 1548 21498
rect 900 21455 1548 21464
rect 162 21412 810 21421
rect 162 21378 810 21412
rect 162 21369 810 21378
rect 900 21326 1548 21335
rect 900 21292 1548 21326
rect 900 21283 1548 21292
rect 162 21240 810 21249
rect 162 21206 810 21240
rect 162 21197 810 21206
rect 900 21154 1548 21163
rect 900 21120 1548 21154
rect 900 21111 1548 21120
rect 162 21068 810 21077
rect 162 21034 810 21068
rect 162 21025 810 21034
rect 900 20982 1548 20991
rect 900 20948 1548 20982
rect 900 20939 1548 20948
rect 162 20896 810 20905
rect 162 20862 810 20896
rect 162 20853 810 20862
rect 900 20810 1548 20819
rect 900 20776 1548 20810
rect 900 20767 1548 20776
rect 162 20724 810 20733
rect 162 20690 810 20724
rect 162 20681 810 20690
rect 900 20638 1548 20647
rect 900 20604 1548 20638
rect 900 20595 1548 20604
rect 162 20552 810 20561
rect 162 20518 810 20552
rect 162 20509 810 20518
rect 900 20466 1548 20475
rect 900 20432 1548 20466
rect 900 20423 1548 20432
rect 162 20380 810 20389
rect 162 20346 810 20380
rect 162 20337 810 20346
rect 900 20294 1548 20303
rect 900 20260 1548 20294
rect 900 20251 1548 20260
rect 162 20208 810 20217
rect 162 20174 810 20208
rect 162 20165 810 20174
rect 900 20122 1548 20131
rect 900 20088 1548 20122
rect 900 20079 1548 20088
rect 162 20036 810 20045
rect 162 20002 810 20036
rect 162 19993 810 20002
rect 900 19950 1548 19959
rect 900 19916 1548 19950
rect 900 19907 1548 19916
rect 162 19864 810 19873
rect 162 19830 810 19864
rect 162 19821 810 19830
rect 900 19778 1548 19787
rect 900 19744 1548 19778
rect 900 19735 1548 19744
rect 162 19692 810 19701
rect 162 19658 810 19692
rect 162 19649 810 19658
rect 900 19606 1548 19615
rect 900 19572 1548 19606
rect 900 19563 1548 19572
rect 162 19520 810 19529
rect 162 19486 810 19520
rect 162 19477 810 19486
rect 900 19434 1548 19443
rect 900 19400 1548 19434
rect 900 19391 1548 19400
rect 162 19348 810 19357
rect 162 19314 810 19348
rect 162 19305 810 19314
rect 900 19262 1548 19271
rect 900 19228 1548 19262
rect 900 19219 1548 19228
rect 162 19176 810 19185
rect 162 19142 810 19176
rect 162 19133 810 19142
rect 900 19090 1548 19099
rect 900 19056 1548 19090
rect 900 19047 1548 19056
rect 162 19004 810 19013
rect 162 18970 810 19004
rect 162 18961 810 18970
rect 900 18918 1548 18927
rect 900 18884 1548 18918
rect 900 18875 1548 18884
rect 162 18832 810 18841
rect 162 18798 810 18832
rect 162 18789 810 18798
rect 900 18746 1548 18755
rect 900 18712 1548 18746
rect 900 18703 1548 18712
rect 162 18660 810 18669
rect 162 18626 810 18660
rect 162 18617 810 18626
rect 900 18574 1548 18583
rect 900 18540 1548 18574
rect 900 18531 1548 18540
rect 162 18488 810 18497
rect 162 18454 810 18488
rect 162 18445 810 18454
rect 900 18402 1548 18411
rect 900 18368 1548 18402
rect 900 18359 1548 18368
rect 162 18316 810 18325
rect 162 18282 810 18316
rect 162 18273 810 18282
rect 900 18230 1548 18239
rect 900 18196 1548 18230
rect 900 18187 1548 18196
rect 162 18144 810 18153
rect 162 18110 810 18144
rect 162 18101 810 18110
rect 900 18058 1548 18067
rect 900 18024 1548 18058
rect 900 18015 1548 18024
rect 162 17972 810 17981
rect 162 17938 810 17972
rect 162 17929 810 17938
rect 900 17886 1548 17895
rect 900 17852 1548 17886
rect 900 17843 1548 17852
rect 162 17800 810 17809
rect 162 17766 810 17800
rect 162 17757 810 17766
rect 900 17714 1548 17723
rect 900 17680 1548 17714
rect 900 17671 1548 17680
rect 162 17628 810 17637
rect 162 17594 810 17628
rect 162 17585 810 17594
rect 900 17542 1548 17551
rect 900 17508 1548 17542
rect 900 17499 1548 17508
rect 162 17456 810 17465
rect 162 17422 810 17456
rect 162 17413 810 17422
rect 900 17370 1548 17379
rect 900 17336 1548 17370
rect 900 17327 1548 17336
rect 162 17284 810 17293
rect 162 17250 810 17284
rect 162 17241 810 17250
rect 900 17198 1548 17207
rect 900 17164 1548 17198
rect 900 17155 1548 17164
rect 162 17112 810 17121
rect 162 17078 810 17112
rect 162 17069 810 17078
rect 900 17026 1548 17035
rect 900 16992 1548 17026
rect 900 16983 1548 16992
rect 162 16940 810 16949
rect 162 16906 810 16940
rect 162 16897 810 16906
rect 900 16854 1548 16863
rect 900 16820 1548 16854
rect 900 16811 1548 16820
rect 162 16768 810 16777
rect 162 16734 810 16768
rect 162 16725 810 16734
rect 900 16682 1548 16691
rect 900 16648 1548 16682
rect 900 16639 1548 16648
rect 162 16596 810 16605
rect 162 16562 810 16596
rect 162 16553 810 16562
rect 900 16510 1548 16519
rect 900 16476 1548 16510
rect 900 16467 1548 16476
rect 162 16424 810 16433
rect 162 16390 810 16424
rect 162 16381 810 16390
rect 900 16338 1548 16347
rect 900 16304 1548 16338
rect 900 16295 1548 16304
rect 162 16252 810 16261
rect 162 16218 810 16252
rect 162 16209 810 16218
rect 900 16166 1548 16175
rect 900 16132 1548 16166
rect 900 16123 1548 16132
rect 162 16080 810 16089
rect 162 16046 810 16080
rect 162 16037 810 16046
rect 900 15994 1548 16003
rect 900 15960 1548 15994
rect 900 15951 1548 15960
rect 162 15908 810 15917
rect 162 15874 810 15908
rect 162 15865 810 15874
rect 900 15822 1548 15831
rect 900 15788 1548 15822
rect 900 15779 1548 15788
rect 162 15736 810 15745
rect 162 15702 810 15736
rect 162 15693 810 15702
rect 900 15650 1548 15659
rect 900 15616 1548 15650
rect 900 15607 1548 15616
rect 162 15564 810 15573
rect 162 15530 810 15564
rect 162 15521 810 15530
rect 900 15478 1548 15487
rect 900 15444 1548 15478
rect 900 15435 1548 15444
rect 162 15392 810 15401
rect 162 15358 810 15392
rect 162 15349 810 15358
rect 900 15306 1548 15315
rect 900 15272 1548 15306
rect 900 15263 1548 15272
rect 162 15220 810 15229
rect 162 15186 810 15220
rect 162 15177 810 15186
rect 900 15134 1548 15143
rect 900 15100 1548 15134
rect 900 15091 1548 15100
rect 162 15048 810 15057
rect 162 15014 810 15048
rect 162 15005 810 15014
rect 900 14962 1548 14971
rect 900 14928 1548 14962
rect 900 14919 1548 14928
rect 162 14876 810 14885
rect 162 14842 810 14876
rect 162 14833 810 14842
rect 900 14790 1548 14799
rect 900 14756 1548 14790
rect 900 14747 1548 14756
rect 162 14704 810 14713
rect 162 14670 810 14704
rect 162 14661 810 14670
rect 900 14618 1548 14627
rect 900 14584 1548 14618
rect 900 14575 1548 14584
rect 162 14532 810 14541
rect 162 14498 810 14532
rect 162 14489 810 14498
rect 900 14446 1548 14455
rect 900 14412 1548 14446
rect 900 14403 1548 14412
rect 162 14360 810 14369
rect 162 14326 810 14360
rect 162 14317 810 14326
rect 900 14274 1548 14283
rect 900 14240 1548 14274
rect 900 14231 1548 14240
rect 162 14188 810 14197
rect 162 14154 810 14188
rect 162 14145 810 14154
rect 900 14102 1548 14111
rect 900 14068 1548 14102
rect 900 14059 1548 14068
rect 162 14016 810 14025
rect 162 13982 810 14016
rect 162 13973 810 13982
rect 900 13930 1548 13939
rect 900 13896 1548 13930
rect 900 13887 1548 13896
rect 162 13844 810 13853
rect 162 13810 810 13844
rect 162 13801 810 13810
rect 900 13758 1548 13767
rect 900 13724 1548 13758
rect 900 13715 1548 13724
rect 162 13672 810 13681
rect 162 13638 810 13672
rect 162 13629 810 13638
rect 900 13586 1548 13595
rect 900 13552 1548 13586
rect 900 13543 1548 13552
rect 162 13500 810 13509
rect 162 13466 810 13500
rect 162 13457 810 13466
rect 900 13414 1548 13423
rect 900 13380 1548 13414
rect 900 13371 1548 13380
rect 162 13328 810 13337
rect 162 13294 810 13328
rect 162 13285 810 13294
rect 900 13242 1548 13251
rect 900 13208 1548 13242
rect 900 13199 1548 13208
rect 162 13156 810 13165
rect 162 13122 810 13156
rect 162 13113 810 13122
rect 900 13070 1548 13079
rect 900 13036 1548 13070
rect 900 13027 1548 13036
rect 162 12984 810 12993
rect 162 12950 810 12984
rect 162 12941 810 12950
rect 900 12898 1548 12907
rect 900 12864 1548 12898
rect 900 12855 1548 12864
rect 162 12812 810 12821
rect 162 12778 810 12812
rect 162 12769 810 12778
rect 900 12726 1548 12735
rect 900 12692 1548 12726
rect 900 12683 1548 12692
rect 162 12640 810 12649
rect 162 12606 810 12640
rect 162 12597 810 12606
rect 900 12554 1548 12563
rect 900 12520 1548 12554
rect 900 12511 1548 12520
rect 162 12468 810 12477
rect 162 12434 810 12468
rect 162 12425 810 12434
rect 900 12382 1548 12391
rect 900 12348 1548 12382
rect 900 12339 1548 12348
rect 162 12296 810 12305
rect 162 12262 810 12296
rect 162 12253 810 12262
rect 900 12210 1548 12219
rect 900 12176 1548 12210
rect 900 12167 1548 12176
rect 162 12124 810 12133
rect 162 12090 810 12124
rect 162 12081 810 12090
rect 900 12038 1548 12047
rect 900 12004 1548 12038
rect 900 11995 1548 12004
rect 162 11952 810 11961
rect 162 11918 810 11952
rect 162 11909 810 11918
rect 900 11866 1548 11875
rect 900 11832 1548 11866
rect 900 11823 1548 11832
rect 162 11780 810 11789
rect 162 11746 810 11780
rect 162 11737 810 11746
rect 900 11694 1548 11703
rect 900 11660 1548 11694
rect 900 11651 1548 11660
rect 162 11608 810 11617
rect 162 11574 810 11608
rect 162 11565 810 11574
rect 900 11522 1548 11531
rect 900 11488 1548 11522
rect 900 11479 1548 11488
rect 162 11436 810 11445
rect 162 11402 810 11436
rect 162 11393 810 11402
rect 900 11350 1548 11359
rect 900 11316 1548 11350
rect 900 11307 1548 11316
rect 162 11264 810 11273
rect 162 11230 810 11264
rect 162 11221 810 11230
rect 900 11178 1548 11187
rect 900 11144 1548 11178
rect 900 11135 1548 11144
rect 162 11092 810 11101
rect 162 11058 810 11092
rect 162 11049 810 11058
rect 900 11006 1548 11015
rect 900 10972 1548 11006
rect 900 10963 1548 10972
rect 162 10920 810 10929
rect 162 10886 810 10920
rect 162 10877 810 10886
rect 900 10834 1548 10843
rect 900 10800 1548 10834
rect 900 10791 1548 10800
rect 162 10748 810 10757
rect 162 10714 810 10748
rect 162 10705 810 10714
rect 900 10662 1548 10671
rect 900 10628 1548 10662
rect 900 10619 1548 10628
rect 162 10576 810 10585
rect 162 10542 810 10576
rect 162 10533 810 10542
rect 900 10490 1548 10499
rect 900 10456 1548 10490
rect 900 10447 1548 10456
rect 162 10404 810 10413
rect 162 10370 810 10404
rect 162 10361 810 10370
rect 900 10318 1548 10327
rect 900 10284 1548 10318
rect 900 10275 1548 10284
rect 162 10232 810 10241
rect 162 10198 810 10232
rect 162 10189 810 10198
rect 900 10146 1548 10155
rect 900 10112 1548 10146
rect 900 10103 1548 10112
rect 162 10060 810 10069
rect 162 10026 810 10060
rect 162 10017 810 10026
rect 900 9974 1548 9983
rect 900 9940 1548 9974
rect 900 9931 1548 9940
rect 162 9888 810 9897
rect 162 9854 810 9888
rect 162 9845 810 9854
rect 900 9802 1548 9811
rect 900 9768 1548 9802
rect 900 9759 1548 9768
rect 162 9716 810 9725
rect 162 9682 810 9716
rect 162 9673 810 9682
rect 900 9630 1548 9639
rect 900 9596 1548 9630
rect 900 9587 1548 9596
rect 162 9544 810 9553
rect 162 9510 810 9544
rect 162 9501 810 9510
rect 900 9458 1548 9467
rect 900 9424 1548 9458
rect 900 9415 1548 9424
rect 162 9372 810 9381
rect 162 9338 810 9372
rect 162 9329 810 9338
rect 900 9286 1548 9295
rect 900 9252 1548 9286
rect 900 9243 1548 9252
rect 162 9200 810 9209
rect 162 9166 810 9200
rect 162 9157 810 9166
rect 900 9114 1548 9123
rect 900 9080 1548 9114
rect 900 9071 1548 9080
rect 162 9028 810 9037
rect 162 8994 810 9028
rect 162 8985 810 8994
rect 900 8942 1548 8951
rect 900 8908 1548 8942
rect 900 8899 1548 8908
rect 162 8856 810 8865
rect 162 8822 810 8856
rect 162 8813 810 8822
rect 900 8770 1548 8779
rect 900 8736 1548 8770
rect 900 8727 1548 8736
rect 162 8684 810 8693
rect 162 8650 810 8684
rect 162 8641 810 8650
rect 900 8598 1548 8607
rect 900 8564 1548 8598
rect 900 8555 1548 8564
rect 162 8512 810 8521
rect 162 8478 810 8512
rect 162 8469 810 8478
rect 900 8426 1548 8435
rect 900 8392 1548 8426
rect 900 8383 1548 8392
rect 162 8340 810 8349
rect 162 8306 810 8340
rect 162 8297 810 8306
rect 900 8254 1548 8263
rect 900 8220 1548 8254
rect 900 8211 1548 8220
rect 162 8168 810 8177
rect 162 8134 810 8168
rect 162 8125 810 8134
rect 900 8082 1548 8091
rect 900 8048 1548 8082
rect 900 8039 1548 8048
rect 162 7996 810 8005
rect 162 7962 810 7996
rect 162 7953 810 7962
rect 900 7910 1548 7919
rect 900 7876 1548 7910
rect 900 7867 1548 7876
rect 162 7824 810 7833
rect 162 7790 810 7824
rect 162 7781 810 7790
rect 900 7738 1548 7747
rect 900 7704 1548 7738
rect 900 7695 1548 7704
rect 162 7652 810 7661
rect 162 7618 810 7652
rect 162 7609 810 7618
rect 900 7566 1548 7575
rect 900 7532 1548 7566
rect 900 7523 1548 7532
rect 162 7480 810 7489
rect 162 7446 810 7480
rect 162 7437 810 7446
rect 900 7394 1548 7403
rect 900 7360 1548 7394
rect 900 7351 1548 7360
rect 162 7308 810 7317
rect 162 7274 810 7308
rect 162 7265 810 7274
rect 900 7222 1548 7231
rect 900 7188 1548 7222
rect 900 7179 1548 7188
rect 162 7136 810 7145
rect 162 7102 810 7136
rect 162 7093 810 7102
rect 900 7050 1548 7059
rect 900 7016 1548 7050
rect 900 7007 1548 7016
rect 162 6964 810 6973
rect 162 6930 810 6964
rect 162 6921 810 6930
rect 900 6878 1548 6887
rect 900 6844 1548 6878
rect 900 6835 1548 6844
rect 162 6792 810 6801
rect 162 6758 810 6792
rect 162 6749 810 6758
rect 900 6706 1548 6715
rect 900 6672 1548 6706
rect 900 6663 1548 6672
rect 162 6620 810 6629
rect 162 6586 810 6620
rect 162 6577 810 6586
rect 900 6534 1548 6543
rect 900 6500 1548 6534
rect 900 6491 1548 6500
rect 162 6448 810 6457
rect 162 6414 810 6448
rect 162 6405 810 6414
rect 900 6362 1548 6371
rect 900 6328 1548 6362
rect 900 6319 1548 6328
rect 162 6276 810 6285
rect 162 6242 810 6276
rect 162 6233 810 6242
rect 900 6190 1548 6199
rect 900 6156 1548 6190
rect 900 6147 1548 6156
rect 162 6104 810 6113
rect 162 6070 810 6104
rect 162 6061 810 6070
rect 900 6018 1548 6027
rect 900 5984 1548 6018
rect 900 5975 1548 5984
rect 162 5932 810 5941
rect 162 5898 810 5932
rect 162 5889 810 5898
rect 900 5846 1548 5855
rect 900 5812 1548 5846
rect 900 5803 1548 5812
rect 162 5760 810 5769
rect 162 5726 810 5760
rect 162 5717 810 5726
rect 900 5674 1548 5683
rect 900 5640 1548 5674
rect 900 5631 1548 5640
rect 162 5588 810 5597
rect 162 5554 810 5588
rect 162 5545 810 5554
rect 900 5502 1548 5511
rect 900 5468 1548 5502
rect 900 5459 1548 5468
rect 162 5416 810 5425
rect 162 5382 810 5416
rect 162 5373 810 5382
rect 900 5330 1548 5339
rect 900 5296 1548 5330
rect 900 5287 1548 5296
rect 162 5244 810 5253
rect 162 5210 810 5244
rect 162 5201 810 5210
rect 900 5158 1548 5167
rect 900 5124 1548 5158
rect 900 5115 1548 5124
rect 162 5072 810 5081
rect 162 5038 810 5072
rect 162 5029 810 5038
rect 900 4986 1548 4995
rect 900 4952 1548 4986
rect 900 4943 1548 4952
rect 162 4900 810 4909
rect 162 4866 810 4900
rect 162 4857 810 4866
rect 900 4814 1548 4823
rect 900 4780 1548 4814
rect 900 4771 1548 4780
rect 162 4728 810 4737
rect 162 4694 810 4728
rect 162 4685 810 4694
rect 900 4642 1548 4651
rect 900 4608 1548 4642
rect 900 4599 1548 4608
rect 162 4556 810 4565
rect 162 4522 810 4556
rect 162 4513 810 4522
rect 900 4470 1548 4479
rect 900 4436 1548 4470
rect 900 4427 1548 4436
rect 162 4384 810 4393
rect 162 4350 810 4384
rect 162 4341 810 4350
rect 900 4298 1548 4307
rect 900 4264 1548 4298
rect 900 4255 1548 4264
rect 162 4212 810 4221
rect 162 4178 810 4212
rect 162 4169 810 4178
rect 900 4126 1548 4135
rect 900 4092 1548 4126
rect 900 4083 1548 4092
rect 162 4040 810 4049
rect 162 4006 810 4040
rect 162 3997 810 4006
rect 900 3954 1548 3963
rect 900 3920 1548 3954
rect 900 3911 1548 3920
rect 162 3868 810 3877
rect 162 3834 810 3868
rect 162 3825 810 3834
rect 900 3782 1548 3791
rect 900 3748 1548 3782
rect 900 3739 1548 3748
rect 162 3696 810 3705
rect 162 3662 810 3696
rect 162 3653 810 3662
rect 900 3610 1548 3619
rect 900 3576 1548 3610
rect 900 3567 1548 3576
rect 162 3524 810 3533
rect 162 3490 810 3524
rect 162 3481 810 3490
rect 900 3438 1548 3447
rect 900 3404 1548 3438
rect 900 3395 1548 3404
rect 162 3352 810 3361
rect 162 3318 810 3352
rect 162 3309 810 3318
rect 900 3266 1548 3275
rect 900 3232 1548 3266
rect 900 3223 1548 3232
rect 162 3180 810 3189
rect 162 3146 810 3180
rect 162 3137 810 3146
rect 900 3094 1548 3103
rect 900 3060 1548 3094
rect 900 3051 1548 3060
rect 162 3008 810 3017
rect 162 2974 810 3008
rect 162 2965 810 2974
rect 900 2922 1548 2931
rect 900 2888 1548 2922
rect 900 2879 1548 2888
rect 162 2836 810 2845
rect 162 2802 810 2836
rect 162 2793 810 2802
rect 900 2750 1548 2759
rect 900 2716 1548 2750
rect 900 2707 1548 2716
rect 162 2664 810 2673
rect 162 2630 810 2664
rect 162 2621 810 2630
rect 900 2578 1548 2587
rect 900 2544 1548 2578
rect 900 2535 1548 2544
rect 162 2492 810 2501
rect 162 2458 810 2492
rect 162 2449 810 2458
rect 900 2406 1548 2415
rect 900 2372 1548 2406
rect 900 2363 1548 2372
rect 162 2320 810 2329
rect 162 2286 810 2320
rect 162 2277 810 2286
rect 900 2234 1548 2243
rect 900 2200 1548 2234
rect 900 2191 1548 2200
rect 162 2148 810 2157
rect 162 2114 810 2148
rect 162 2105 810 2114
rect 900 2062 1548 2071
rect 900 2028 1548 2062
rect 900 2019 1548 2028
rect 162 1976 810 1985
rect 162 1942 810 1976
rect 162 1933 810 1942
rect 900 1890 1548 1899
rect 900 1856 1548 1890
rect 900 1847 1548 1856
rect 162 1804 810 1813
rect 162 1770 810 1804
rect 162 1761 810 1770
rect 900 1718 1548 1727
rect 900 1684 1548 1718
rect 900 1675 1548 1684
rect 162 1632 810 1641
rect 162 1598 810 1632
rect 162 1589 810 1598
rect 900 1546 1548 1555
rect 900 1512 1548 1546
rect 900 1503 1548 1512
rect 162 1460 810 1469
rect 162 1426 810 1460
rect 162 1417 810 1426
rect 900 1374 1548 1383
rect 900 1340 1548 1374
rect 900 1331 1548 1340
rect 162 1288 810 1297
rect 162 1254 810 1288
rect 162 1245 810 1254
rect 900 1202 1548 1211
rect 900 1168 1548 1202
rect 900 1159 1548 1168
rect 162 1116 810 1125
rect 162 1082 810 1116
rect 162 1073 810 1082
rect 900 1030 1548 1039
rect 900 996 1548 1030
rect 900 987 1548 996
rect 162 944 810 953
rect 162 910 810 944
rect 162 901 810 910
rect 900 858 1548 867
rect 900 824 1548 858
rect 900 815 1548 824
rect 162 772 810 781
rect 162 738 810 772
rect 162 729 810 738
rect 900 686 1548 695
rect 900 652 1548 686
rect 900 643 1548 652
rect 162 600 810 609
rect 162 566 810 600
rect 162 557 810 566
rect 900 514 1548 523
rect 900 480 1548 514
rect 900 471 1548 480
rect 162 428 810 437
rect 162 394 810 428
rect 162 385 810 394
rect 900 342 1548 351
rect 900 308 1548 342
rect 900 299 1548 308
rect 162 256 810 265
rect 162 222 810 256
rect 162 213 810 222
rect 1618 179 1628 43815
rect 1628 179 1662 43815
rect 1662 179 1672 43815
rect 900 170 1548 179
rect 900 136 1548 170
rect 1618 169 1672 179
rect 900 127 1548 136
<< metal2 >>
rect 156 43781 816 43867
rect 156 43729 162 43781
rect 810 43729 816 43781
rect 156 43609 816 43729
rect 156 43557 162 43609
rect 810 43557 816 43609
rect 156 43437 816 43557
rect 156 43385 162 43437
rect 810 43385 816 43437
rect 156 43265 816 43385
rect 156 43213 162 43265
rect 810 43213 816 43265
rect 156 43093 816 43213
rect 156 43041 162 43093
rect 810 43041 816 43093
rect 156 42921 816 43041
rect 156 42869 162 42921
rect 810 42869 816 42921
rect 156 42749 816 42869
rect 156 42697 162 42749
rect 810 42697 816 42749
rect 156 42577 816 42697
rect 156 42525 162 42577
rect 810 42525 816 42577
rect 156 42405 816 42525
rect 156 42353 162 42405
rect 810 42353 816 42405
rect 156 42233 816 42353
rect 156 42181 162 42233
rect 810 42181 816 42233
rect 156 42061 816 42181
rect 156 42009 162 42061
rect 810 42009 816 42061
rect 156 41889 816 42009
rect 156 41837 162 41889
rect 810 41837 816 41889
rect 156 41717 816 41837
rect 156 41665 162 41717
rect 810 41665 816 41717
rect 156 41545 816 41665
rect 156 41493 162 41545
rect 810 41493 816 41545
rect 156 41373 816 41493
rect 156 41321 162 41373
rect 810 41321 816 41373
rect 156 41201 816 41321
rect 156 41149 162 41201
rect 810 41149 816 41201
rect 156 41029 816 41149
rect 156 40977 162 41029
rect 810 40977 816 41029
rect 156 40857 816 40977
rect 156 40805 162 40857
rect 810 40805 816 40857
rect 156 40685 816 40805
rect 156 40633 162 40685
rect 810 40633 816 40685
rect 156 40513 816 40633
rect 156 40461 162 40513
rect 810 40461 816 40513
rect 156 40341 816 40461
rect 156 40289 162 40341
rect 810 40289 816 40341
rect 156 40169 816 40289
rect 156 40117 162 40169
rect 810 40117 816 40169
rect 156 39997 816 40117
rect 156 39945 162 39997
rect 810 39945 816 39997
rect 156 39825 816 39945
rect 156 39773 162 39825
rect 810 39773 816 39825
rect 156 39653 816 39773
rect 156 39601 162 39653
rect 810 39601 816 39653
rect 156 39481 816 39601
rect 156 39429 162 39481
rect 810 39429 816 39481
rect 156 39309 816 39429
rect 156 39257 162 39309
rect 810 39257 816 39309
rect 156 39137 816 39257
rect 156 39085 162 39137
rect 810 39085 816 39137
rect 156 38965 816 39085
rect 156 38913 162 38965
rect 810 38913 816 38965
rect 156 38793 816 38913
rect 156 38741 162 38793
rect 810 38741 816 38793
rect 156 38621 816 38741
rect 156 38569 162 38621
rect 810 38569 816 38621
rect 156 38449 816 38569
rect 156 38397 162 38449
rect 810 38397 816 38449
rect 156 38277 816 38397
rect 156 38225 162 38277
rect 810 38225 816 38277
rect 156 38105 816 38225
rect 156 38053 162 38105
rect 810 38053 816 38105
rect 156 37933 816 38053
rect 156 37881 162 37933
rect 810 37881 816 37933
rect 156 37761 816 37881
rect 156 37709 162 37761
rect 810 37709 816 37761
rect 156 37589 816 37709
rect 156 37537 162 37589
rect 810 37537 816 37589
rect 156 37417 816 37537
rect 156 37365 162 37417
rect 810 37365 816 37417
rect 156 37245 816 37365
rect 156 37193 162 37245
rect 810 37193 816 37245
rect 156 37073 816 37193
rect 156 37021 162 37073
rect 810 37021 816 37073
rect 156 36901 816 37021
rect 156 36849 162 36901
rect 810 36849 816 36901
rect 156 36729 816 36849
rect 156 36677 162 36729
rect 810 36677 816 36729
rect 156 36557 816 36677
rect 156 36505 162 36557
rect 810 36505 816 36557
rect 156 36385 816 36505
rect 156 36333 162 36385
rect 810 36333 816 36385
rect 156 36213 816 36333
rect 156 36161 162 36213
rect 810 36161 816 36213
rect 156 36041 816 36161
rect 156 35989 162 36041
rect 810 35989 816 36041
rect 156 35869 816 35989
rect 156 35817 162 35869
rect 810 35817 816 35869
rect 156 35697 816 35817
rect 156 35645 162 35697
rect 810 35645 816 35697
rect 156 35525 816 35645
rect 156 35473 162 35525
rect 810 35473 816 35525
rect 156 35353 816 35473
rect 156 35301 162 35353
rect 810 35301 816 35353
rect 156 35181 816 35301
rect 156 35129 162 35181
rect 810 35129 816 35181
rect 156 35009 816 35129
rect 156 34957 162 35009
rect 810 34957 816 35009
rect 156 34837 816 34957
rect 156 34785 162 34837
rect 810 34785 816 34837
rect 156 34665 816 34785
rect 156 34613 162 34665
rect 810 34613 816 34665
rect 156 34493 816 34613
rect 156 34441 162 34493
rect 810 34441 816 34493
rect 156 34321 816 34441
rect 156 34269 162 34321
rect 810 34269 816 34321
rect 156 34149 816 34269
rect 156 34097 162 34149
rect 810 34097 816 34149
rect 156 33977 816 34097
rect 156 33925 162 33977
rect 810 33925 816 33977
rect 156 33805 816 33925
rect 156 33753 162 33805
rect 810 33753 816 33805
rect 156 33633 816 33753
rect 156 33581 162 33633
rect 810 33581 816 33633
rect 156 33461 816 33581
rect 156 33409 162 33461
rect 810 33409 816 33461
rect 156 33289 816 33409
rect 156 33237 162 33289
rect 810 33237 816 33289
rect 156 33117 816 33237
rect 156 33065 162 33117
rect 810 33065 816 33117
rect 156 32945 816 33065
rect 156 32893 162 32945
rect 810 32893 816 32945
rect 156 32773 816 32893
rect 156 32721 162 32773
rect 810 32721 816 32773
rect 156 32601 816 32721
rect 156 32549 162 32601
rect 810 32549 816 32601
rect 156 32429 816 32549
rect 156 32377 162 32429
rect 810 32377 816 32429
rect 156 32257 816 32377
rect 156 32205 162 32257
rect 810 32205 816 32257
rect 156 32085 816 32205
rect 156 32033 162 32085
rect 810 32033 816 32085
rect 156 31913 816 32033
rect 156 31861 162 31913
rect 810 31861 816 31913
rect 156 31741 816 31861
rect 156 31689 162 31741
rect 810 31689 816 31741
rect 156 31569 816 31689
rect 156 31517 162 31569
rect 810 31517 816 31569
rect 156 31397 816 31517
rect 156 31345 162 31397
rect 810 31345 816 31397
rect 156 31225 816 31345
rect 156 31173 162 31225
rect 810 31173 816 31225
rect 156 31053 816 31173
rect 156 31001 162 31053
rect 810 31001 816 31053
rect 156 30881 816 31001
rect 156 30829 162 30881
rect 810 30829 816 30881
rect 156 30709 816 30829
rect 156 30657 162 30709
rect 810 30657 816 30709
rect 156 30537 816 30657
rect 156 30485 162 30537
rect 810 30485 816 30537
rect 156 30365 816 30485
rect 156 30313 162 30365
rect 810 30313 816 30365
rect 156 30193 816 30313
rect 156 30141 162 30193
rect 810 30141 816 30193
rect 156 30021 816 30141
rect 156 29969 162 30021
rect 810 29969 816 30021
rect 156 29849 816 29969
rect 156 29797 162 29849
rect 810 29797 816 29849
rect 156 29677 816 29797
rect 156 29625 162 29677
rect 810 29625 816 29677
rect 156 29505 816 29625
rect 156 29453 162 29505
rect 810 29453 816 29505
rect 156 29333 816 29453
rect 156 29281 162 29333
rect 810 29281 816 29333
rect 156 29161 816 29281
rect 156 29109 162 29161
rect 810 29109 816 29161
rect 156 28989 816 29109
rect 156 28937 162 28989
rect 810 28937 816 28989
rect 156 28817 816 28937
rect 156 28765 162 28817
rect 810 28765 816 28817
rect 156 28645 816 28765
rect 156 28593 162 28645
rect 810 28593 816 28645
rect 156 28473 816 28593
rect 156 28421 162 28473
rect 810 28421 816 28473
rect 156 28301 816 28421
rect 156 28249 162 28301
rect 810 28249 816 28301
rect 156 28129 816 28249
rect 156 28077 162 28129
rect 810 28077 816 28129
rect 156 27957 816 28077
rect 156 27905 162 27957
rect 810 27905 816 27957
rect 156 27785 816 27905
rect 156 27733 162 27785
rect 810 27733 816 27785
rect 156 27613 816 27733
rect 156 27561 162 27613
rect 810 27561 816 27613
rect 156 27441 816 27561
rect 156 27389 162 27441
rect 810 27389 816 27441
rect 156 27269 816 27389
rect 156 27217 162 27269
rect 810 27217 816 27269
rect 156 27097 816 27217
rect 156 27045 162 27097
rect 810 27045 816 27097
rect 156 26925 816 27045
rect 156 26873 162 26925
rect 810 26873 816 26925
rect 156 26753 816 26873
rect 156 26701 162 26753
rect 810 26701 816 26753
rect 156 26581 816 26701
rect 156 26529 162 26581
rect 810 26529 816 26581
rect 156 26409 816 26529
rect 156 26357 162 26409
rect 810 26357 816 26409
rect 156 26237 816 26357
rect 156 26185 162 26237
rect 810 26185 816 26237
rect 156 26065 816 26185
rect 156 26013 162 26065
rect 810 26013 816 26065
rect 156 25893 816 26013
rect 156 25841 162 25893
rect 810 25841 816 25893
rect 156 25721 816 25841
rect 156 25669 162 25721
rect 810 25669 816 25721
rect 156 25549 816 25669
rect 156 25497 162 25549
rect 810 25497 816 25549
rect 156 25377 816 25497
rect 156 25325 162 25377
rect 810 25325 816 25377
rect 156 25205 816 25325
rect 156 25153 162 25205
rect 810 25153 816 25205
rect 156 25033 816 25153
rect 156 24981 162 25033
rect 810 24981 816 25033
rect 156 24861 816 24981
rect 156 24809 162 24861
rect 810 24809 816 24861
rect 156 24689 816 24809
rect 156 24637 162 24689
rect 810 24637 816 24689
rect 156 24517 816 24637
rect 156 24465 162 24517
rect 810 24465 816 24517
rect 156 24345 816 24465
rect 156 24293 162 24345
rect 810 24293 816 24345
rect 156 24173 816 24293
rect 156 24121 162 24173
rect 810 24121 816 24173
rect 156 24001 816 24121
rect 156 23949 162 24001
rect 810 23949 816 24001
rect 156 23829 816 23949
rect 156 23777 162 23829
rect 810 23777 816 23829
rect 156 23657 816 23777
rect 156 23605 162 23657
rect 810 23605 816 23657
rect 156 23485 816 23605
rect 156 23433 162 23485
rect 810 23433 816 23485
rect 156 23313 816 23433
rect 156 23261 162 23313
rect 810 23261 816 23313
rect 156 23141 816 23261
rect 156 23089 162 23141
rect 810 23089 816 23141
rect 156 22969 816 23089
rect 156 22917 162 22969
rect 810 22917 816 22969
rect 156 22797 816 22917
rect 156 22745 162 22797
rect 810 22745 816 22797
rect 156 22625 816 22745
rect 156 22573 162 22625
rect 810 22573 816 22625
rect 156 22453 816 22573
rect 156 22401 162 22453
rect 810 22401 816 22453
rect 156 22281 816 22401
rect 156 22229 162 22281
rect 810 22229 816 22281
rect 156 22109 816 22229
rect 156 22057 162 22109
rect 810 22057 816 22109
rect 156 21937 816 22057
rect 156 21885 162 21937
rect 810 21885 816 21937
rect 156 21765 816 21885
rect 156 21713 162 21765
rect 810 21713 816 21765
rect 156 21593 816 21713
rect 156 21541 162 21593
rect 810 21541 816 21593
rect 156 21421 816 21541
rect 156 21369 162 21421
rect 810 21369 816 21421
rect 156 21249 816 21369
rect 156 21197 162 21249
rect 810 21197 816 21249
rect 156 21077 816 21197
rect 156 21025 162 21077
rect 810 21025 816 21077
rect 156 20905 816 21025
rect 156 20853 162 20905
rect 810 20853 816 20905
rect 156 20733 816 20853
rect 156 20681 162 20733
rect 810 20681 816 20733
rect 156 20561 816 20681
rect 156 20509 162 20561
rect 810 20509 816 20561
rect 156 20389 816 20509
rect 156 20337 162 20389
rect 810 20337 816 20389
rect 156 20217 816 20337
rect 156 20165 162 20217
rect 810 20165 816 20217
rect 156 20045 816 20165
rect 156 19993 162 20045
rect 810 19993 816 20045
rect 156 19873 816 19993
rect 156 19821 162 19873
rect 810 19821 816 19873
rect 156 19701 816 19821
rect 156 19649 162 19701
rect 810 19649 816 19701
rect 156 19529 816 19649
rect 156 19477 162 19529
rect 810 19477 816 19529
rect 156 19357 816 19477
rect 156 19305 162 19357
rect 810 19305 816 19357
rect 156 19185 816 19305
rect 156 19133 162 19185
rect 810 19133 816 19185
rect 156 19013 816 19133
rect 156 18961 162 19013
rect 810 18961 816 19013
rect 156 18841 816 18961
rect 156 18789 162 18841
rect 810 18789 816 18841
rect 156 18669 816 18789
rect 156 18617 162 18669
rect 810 18617 816 18669
rect 156 18497 816 18617
rect 156 18445 162 18497
rect 810 18445 816 18497
rect 156 18325 816 18445
rect 156 18273 162 18325
rect 810 18273 816 18325
rect 156 18153 816 18273
rect 156 18101 162 18153
rect 810 18101 816 18153
rect 156 17981 816 18101
rect 156 17929 162 17981
rect 810 17929 816 17981
rect 156 17809 816 17929
rect 156 17757 162 17809
rect 810 17757 816 17809
rect 156 17637 816 17757
rect 156 17585 162 17637
rect 810 17585 816 17637
rect 156 17465 816 17585
rect 156 17413 162 17465
rect 810 17413 816 17465
rect 156 17293 816 17413
rect 156 17241 162 17293
rect 810 17241 816 17293
rect 156 17121 816 17241
rect 156 17069 162 17121
rect 810 17069 816 17121
rect 156 16949 816 17069
rect 156 16897 162 16949
rect 810 16897 816 16949
rect 156 16777 816 16897
rect 156 16725 162 16777
rect 810 16725 816 16777
rect 156 16605 816 16725
rect 156 16553 162 16605
rect 810 16553 816 16605
rect 156 16433 816 16553
rect 156 16381 162 16433
rect 810 16381 816 16433
rect 156 16261 816 16381
rect 156 16209 162 16261
rect 810 16209 816 16261
rect 156 16089 816 16209
rect 156 16037 162 16089
rect 810 16037 816 16089
rect 156 15917 816 16037
rect 156 15865 162 15917
rect 810 15865 816 15917
rect 156 15745 816 15865
rect 156 15693 162 15745
rect 810 15693 816 15745
rect 156 15573 816 15693
rect 156 15521 162 15573
rect 810 15521 816 15573
rect 156 15401 816 15521
rect 156 15349 162 15401
rect 810 15349 816 15401
rect 156 15229 816 15349
rect 156 15177 162 15229
rect 810 15177 816 15229
rect 156 15057 816 15177
rect 156 15005 162 15057
rect 810 15005 816 15057
rect 156 14885 816 15005
rect 156 14833 162 14885
rect 810 14833 816 14885
rect 156 14713 816 14833
rect 156 14661 162 14713
rect 810 14661 816 14713
rect 156 14541 816 14661
rect 156 14489 162 14541
rect 810 14489 816 14541
rect 156 14369 816 14489
rect 156 14317 162 14369
rect 810 14317 816 14369
rect 156 14197 816 14317
rect 156 14145 162 14197
rect 810 14145 816 14197
rect 156 14025 816 14145
rect 156 13973 162 14025
rect 810 13973 816 14025
rect 156 13853 816 13973
rect 156 13801 162 13853
rect 810 13801 816 13853
rect 156 13681 816 13801
rect 156 13629 162 13681
rect 810 13629 816 13681
rect 156 13509 816 13629
rect 156 13457 162 13509
rect 810 13457 816 13509
rect 156 13337 816 13457
rect 156 13285 162 13337
rect 810 13285 816 13337
rect 156 13165 816 13285
rect 156 13113 162 13165
rect 810 13113 816 13165
rect 156 12993 816 13113
rect 156 12941 162 12993
rect 810 12941 816 12993
rect 156 12821 816 12941
rect 156 12769 162 12821
rect 810 12769 816 12821
rect 156 12649 816 12769
rect 156 12597 162 12649
rect 810 12597 816 12649
rect 156 12477 816 12597
rect 156 12425 162 12477
rect 810 12425 816 12477
rect 156 12305 816 12425
rect 156 12253 162 12305
rect 810 12253 816 12305
rect 156 12133 816 12253
rect 156 12081 162 12133
rect 810 12081 816 12133
rect 156 11961 816 12081
rect 156 11909 162 11961
rect 810 11909 816 11961
rect 156 11789 816 11909
rect 156 11737 162 11789
rect 810 11737 816 11789
rect 156 11617 816 11737
rect 156 11565 162 11617
rect 810 11565 816 11617
rect 156 11445 816 11565
rect 156 11393 162 11445
rect 810 11393 816 11445
rect 156 11273 816 11393
rect 156 11221 162 11273
rect 810 11221 816 11273
rect 156 11101 816 11221
rect 156 11049 162 11101
rect 810 11049 816 11101
rect 156 10929 816 11049
rect 156 10877 162 10929
rect 810 10877 816 10929
rect 156 10757 816 10877
rect 156 10705 162 10757
rect 810 10705 816 10757
rect 156 10585 816 10705
rect 156 10533 162 10585
rect 810 10533 816 10585
rect 156 10413 816 10533
rect 156 10361 162 10413
rect 810 10361 816 10413
rect 156 10241 816 10361
rect 156 10189 162 10241
rect 810 10189 816 10241
rect 156 10069 816 10189
rect 156 10017 162 10069
rect 810 10017 816 10069
rect 156 9897 816 10017
rect 156 9845 162 9897
rect 810 9845 816 9897
rect 156 9725 816 9845
rect 156 9673 162 9725
rect 810 9673 816 9725
rect 156 9553 816 9673
rect 156 9501 162 9553
rect 810 9501 816 9553
rect 156 9381 816 9501
rect 156 9329 162 9381
rect 810 9329 816 9381
rect 156 9209 816 9329
rect 156 9157 162 9209
rect 810 9157 816 9209
rect 156 9037 816 9157
rect 156 8985 162 9037
rect 810 8985 816 9037
rect 156 8865 816 8985
rect 156 8813 162 8865
rect 810 8813 816 8865
rect 156 8693 816 8813
rect 156 8641 162 8693
rect 810 8641 816 8693
rect 156 8521 816 8641
rect 156 8469 162 8521
rect 810 8469 816 8521
rect 156 8349 816 8469
rect 156 8297 162 8349
rect 810 8297 816 8349
rect 156 8177 816 8297
rect 156 8125 162 8177
rect 810 8125 816 8177
rect 156 8005 816 8125
rect 156 7953 162 8005
rect 810 7953 816 8005
rect 156 7833 816 7953
rect 156 7781 162 7833
rect 810 7781 816 7833
rect 156 7661 816 7781
rect 156 7609 162 7661
rect 810 7609 816 7661
rect 156 7489 816 7609
rect 156 7437 162 7489
rect 810 7437 816 7489
rect 156 7317 816 7437
rect 156 7265 162 7317
rect 810 7265 816 7317
rect 156 7145 816 7265
rect 156 7093 162 7145
rect 810 7093 816 7145
rect 156 6973 816 7093
rect 156 6921 162 6973
rect 810 6921 816 6973
rect 156 6801 816 6921
rect 156 6749 162 6801
rect 810 6749 816 6801
rect 156 6629 816 6749
rect 156 6577 162 6629
rect 810 6577 816 6629
rect 156 6457 816 6577
rect 156 6405 162 6457
rect 810 6405 816 6457
rect 156 6285 816 6405
rect 156 6233 162 6285
rect 810 6233 816 6285
rect 156 6113 816 6233
rect 156 6061 162 6113
rect 810 6061 816 6113
rect 156 5941 816 6061
rect 156 5889 162 5941
rect 810 5889 816 5941
rect 156 5769 816 5889
rect 156 5717 162 5769
rect 810 5717 816 5769
rect 156 5597 816 5717
rect 156 5545 162 5597
rect 810 5545 816 5597
rect 156 5425 816 5545
rect 156 5373 162 5425
rect 810 5373 816 5425
rect 156 5253 816 5373
rect 156 5201 162 5253
rect 810 5201 816 5253
rect 156 5081 816 5201
rect 156 5029 162 5081
rect 810 5029 816 5081
rect 156 4909 816 5029
rect 156 4857 162 4909
rect 810 4857 816 4909
rect 156 4737 816 4857
rect 156 4685 162 4737
rect 810 4685 816 4737
rect 156 4565 816 4685
rect 156 4513 162 4565
rect 810 4513 816 4565
rect 156 4393 816 4513
rect 156 4341 162 4393
rect 810 4341 816 4393
rect 156 4221 816 4341
rect 156 4169 162 4221
rect 810 4169 816 4221
rect 156 4049 816 4169
rect 156 3997 162 4049
rect 810 3997 816 4049
rect 156 3877 816 3997
rect 156 3825 162 3877
rect 810 3825 816 3877
rect 156 3705 816 3825
rect 156 3653 162 3705
rect 810 3653 816 3705
rect 156 3533 816 3653
rect 156 3481 162 3533
rect 810 3481 816 3533
rect 156 3361 816 3481
rect 156 3309 162 3361
rect 810 3309 816 3361
rect 156 3189 816 3309
rect 156 3137 162 3189
rect 810 3137 816 3189
rect 156 3017 816 3137
rect 156 2965 162 3017
rect 810 2965 816 3017
rect 156 2845 816 2965
rect 156 2793 162 2845
rect 810 2793 816 2845
rect 156 2673 816 2793
rect 156 2621 162 2673
rect 810 2621 816 2673
rect 156 2501 816 2621
rect 156 2449 162 2501
rect 810 2449 816 2501
rect 156 2329 816 2449
rect 156 2277 162 2329
rect 810 2277 816 2329
rect 156 2157 816 2277
rect 156 2105 162 2157
rect 810 2105 816 2157
rect 156 1985 816 2105
rect 156 1933 162 1985
rect 810 1933 816 1985
rect 156 1813 816 1933
rect 156 1761 162 1813
rect 810 1761 816 1813
rect 156 1641 816 1761
rect 156 1589 162 1641
rect 810 1589 816 1641
rect 156 1469 816 1589
rect 156 1417 162 1469
rect 810 1417 816 1469
rect 156 1297 816 1417
rect 156 1245 162 1297
rect 810 1245 816 1297
rect 156 1125 816 1245
rect 156 1073 162 1125
rect 810 1073 816 1125
rect 156 953 816 1073
rect 156 901 162 953
rect 810 901 816 953
rect 156 781 816 901
rect 156 729 162 781
rect 810 729 816 781
rect 156 609 816 729
rect 156 557 162 609
rect 810 557 816 609
rect 156 437 816 557
rect 156 385 162 437
rect 810 385 816 437
rect 156 265 816 385
rect 156 213 162 265
rect 810 213 816 265
rect 156 127 816 213
rect 894 43815 900 43867
rect 1548 43815 1554 43867
rect 894 43695 1554 43815
rect 894 43643 900 43695
rect 1548 43643 1554 43695
rect 894 43523 1554 43643
rect 894 43471 900 43523
rect 1548 43471 1554 43523
rect 894 43351 1554 43471
rect 894 43299 900 43351
rect 1548 43299 1554 43351
rect 894 43179 1554 43299
rect 894 43127 900 43179
rect 1548 43127 1554 43179
rect 894 43007 1554 43127
rect 894 42955 900 43007
rect 1548 42955 1554 43007
rect 894 42835 1554 42955
rect 894 42783 900 42835
rect 1548 42783 1554 42835
rect 894 42663 1554 42783
rect 894 42611 900 42663
rect 1548 42611 1554 42663
rect 894 42491 1554 42611
rect 894 42439 900 42491
rect 1548 42439 1554 42491
rect 894 42319 1554 42439
rect 894 42267 900 42319
rect 1548 42267 1554 42319
rect 894 42147 1554 42267
rect 894 42095 900 42147
rect 1548 42095 1554 42147
rect 894 41975 1554 42095
rect 894 41923 900 41975
rect 1548 41923 1554 41975
rect 894 41803 1554 41923
rect 894 41751 900 41803
rect 1548 41751 1554 41803
rect 894 41631 1554 41751
rect 894 41579 900 41631
rect 1548 41579 1554 41631
rect 894 41459 1554 41579
rect 894 41407 900 41459
rect 1548 41407 1554 41459
rect 894 41287 1554 41407
rect 894 41235 900 41287
rect 1548 41235 1554 41287
rect 894 41115 1554 41235
rect 894 41063 900 41115
rect 1548 41063 1554 41115
rect 894 40943 1554 41063
rect 894 40891 900 40943
rect 1548 40891 1554 40943
rect 894 40771 1554 40891
rect 894 40719 900 40771
rect 1548 40719 1554 40771
rect 894 40599 1554 40719
rect 894 40547 900 40599
rect 1548 40547 1554 40599
rect 894 40427 1554 40547
rect 894 40375 900 40427
rect 1548 40375 1554 40427
rect 894 40255 1554 40375
rect 894 40203 900 40255
rect 1548 40203 1554 40255
rect 894 40083 1554 40203
rect 894 40031 900 40083
rect 1548 40031 1554 40083
rect 894 39911 1554 40031
rect 894 39859 900 39911
rect 1548 39859 1554 39911
rect 894 39739 1554 39859
rect 894 39687 900 39739
rect 1548 39687 1554 39739
rect 894 39567 1554 39687
rect 894 39515 900 39567
rect 1548 39515 1554 39567
rect 894 39395 1554 39515
rect 894 39343 900 39395
rect 1548 39343 1554 39395
rect 894 39223 1554 39343
rect 894 39171 900 39223
rect 1548 39171 1554 39223
rect 894 39051 1554 39171
rect 894 38999 900 39051
rect 1548 38999 1554 39051
rect 894 38879 1554 38999
rect 894 38827 900 38879
rect 1548 38827 1554 38879
rect 894 38707 1554 38827
rect 894 38655 900 38707
rect 1548 38655 1554 38707
rect 894 38535 1554 38655
rect 894 38483 900 38535
rect 1548 38483 1554 38535
rect 894 38363 1554 38483
rect 894 38311 900 38363
rect 1548 38311 1554 38363
rect 894 38191 1554 38311
rect 894 38139 900 38191
rect 1548 38139 1554 38191
rect 894 38019 1554 38139
rect 894 37967 900 38019
rect 1548 37967 1554 38019
rect 894 37847 1554 37967
rect 894 37795 900 37847
rect 1548 37795 1554 37847
rect 894 37675 1554 37795
rect 894 37623 900 37675
rect 1548 37623 1554 37675
rect 894 37503 1554 37623
rect 894 37451 900 37503
rect 1548 37451 1554 37503
rect 894 37331 1554 37451
rect 894 37279 900 37331
rect 1548 37279 1554 37331
rect 894 37159 1554 37279
rect 894 37107 900 37159
rect 1548 37107 1554 37159
rect 894 36987 1554 37107
rect 894 36935 900 36987
rect 1548 36935 1554 36987
rect 894 36815 1554 36935
rect 894 36763 900 36815
rect 1548 36763 1554 36815
rect 894 36643 1554 36763
rect 894 36591 900 36643
rect 1548 36591 1554 36643
rect 894 36471 1554 36591
rect 894 36419 900 36471
rect 1548 36419 1554 36471
rect 894 36299 1554 36419
rect 894 36247 900 36299
rect 1548 36247 1554 36299
rect 894 36127 1554 36247
rect 894 36075 900 36127
rect 1548 36075 1554 36127
rect 894 35955 1554 36075
rect 894 35903 900 35955
rect 1548 35903 1554 35955
rect 894 35783 1554 35903
rect 894 35731 900 35783
rect 1548 35731 1554 35783
rect 894 35611 1554 35731
rect 894 35559 900 35611
rect 1548 35559 1554 35611
rect 894 35439 1554 35559
rect 894 35387 900 35439
rect 1548 35387 1554 35439
rect 894 35267 1554 35387
rect 894 35215 900 35267
rect 1548 35215 1554 35267
rect 894 35095 1554 35215
rect 894 35043 900 35095
rect 1548 35043 1554 35095
rect 894 34923 1554 35043
rect 894 34871 900 34923
rect 1548 34871 1554 34923
rect 894 34751 1554 34871
rect 894 34699 900 34751
rect 1548 34699 1554 34751
rect 894 34579 1554 34699
rect 894 34527 900 34579
rect 1548 34527 1554 34579
rect 894 34407 1554 34527
rect 894 34355 900 34407
rect 1548 34355 1554 34407
rect 894 34235 1554 34355
rect 894 34183 900 34235
rect 1548 34183 1554 34235
rect 894 34063 1554 34183
rect 894 34011 900 34063
rect 1548 34011 1554 34063
rect 894 33891 1554 34011
rect 894 33839 900 33891
rect 1548 33839 1554 33891
rect 894 33719 1554 33839
rect 894 33667 900 33719
rect 1548 33667 1554 33719
rect 894 33547 1554 33667
rect 894 33495 900 33547
rect 1548 33495 1554 33547
rect 894 33375 1554 33495
rect 894 33323 900 33375
rect 1548 33323 1554 33375
rect 894 33203 1554 33323
rect 894 33151 900 33203
rect 1548 33151 1554 33203
rect 894 33031 1554 33151
rect 894 32979 900 33031
rect 1548 32979 1554 33031
rect 894 32859 1554 32979
rect 894 32807 900 32859
rect 1548 32807 1554 32859
rect 894 32687 1554 32807
rect 894 32635 900 32687
rect 1548 32635 1554 32687
rect 894 32515 1554 32635
rect 894 32463 900 32515
rect 1548 32463 1554 32515
rect 894 32343 1554 32463
rect 894 32291 900 32343
rect 1548 32291 1554 32343
rect 894 32171 1554 32291
rect 894 32119 900 32171
rect 1548 32119 1554 32171
rect 894 31999 1554 32119
rect 894 31947 900 31999
rect 1548 31947 1554 31999
rect 894 31827 1554 31947
rect 894 31775 900 31827
rect 1548 31775 1554 31827
rect 894 31655 1554 31775
rect 894 31603 900 31655
rect 1548 31603 1554 31655
rect 894 31483 1554 31603
rect 894 31431 900 31483
rect 1548 31431 1554 31483
rect 894 31311 1554 31431
rect 894 31259 900 31311
rect 1548 31259 1554 31311
rect 894 31139 1554 31259
rect 894 31087 900 31139
rect 1548 31087 1554 31139
rect 894 30967 1554 31087
rect 894 30915 900 30967
rect 1548 30915 1554 30967
rect 894 30795 1554 30915
rect 894 30743 900 30795
rect 1548 30743 1554 30795
rect 894 30623 1554 30743
rect 894 30571 900 30623
rect 1548 30571 1554 30623
rect 894 30451 1554 30571
rect 894 30399 900 30451
rect 1548 30399 1554 30451
rect 894 30279 1554 30399
rect 894 30227 900 30279
rect 1548 30227 1554 30279
rect 894 30107 1554 30227
rect 894 30055 900 30107
rect 1548 30055 1554 30107
rect 894 29935 1554 30055
rect 894 29883 900 29935
rect 1548 29883 1554 29935
rect 894 29763 1554 29883
rect 894 29711 900 29763
rect 1548 29711 1554 29763
rect 894 29591 1554 29711
rect 894 29539 900 29591
rect 1548 29539 1554 29591
rect 894 29419 1554 29539
rect 894 29367 900 29419
rect 1548 29367 1554 29419
rect 894 29247 1554 29367
rect 894 29195 900 29247
rect 1548 29195 1554 29247
rect 894 29075 1554 29195
rect 894 29023 900 29075
rect 1548 29023 1554 29075
rect 894 28903 1554 29023
rect 894 28851 900 28903
rect 1548 28851 1554 28903
rect 894 28731 1554 28851
rect 894 28679 900 28731
rect 1548 28679 1554 28731
rect 894 28559 1554 28679
rect 894 28507 900 28559
rect 1548 28507 1554 28559
rect 894 28387 1554 28507
rect 894 28335 900 28387
rect 1548 28335 1554 28387
rect 894 28215 1554 28335
rect 894 28163 900 28215
rect 1548 28163 1554 28215
rect 894 28043 1554 28163
rect 894 27991 900 28043
rect 1548 27991 1554 28043
rect 894 27871 1554 27991
rect 894 27819 900 27871
rect 1548 27819 1554 27871
rect 894 27699 1554 27819
rect 894 27647 900 27699
rect 1548 27647 1554 27699
rect 894 27527 1554 27647
rect 894 27475 900 27527
rect 1548 27475 1554 27527
rect 894 27355 1554 27475
rect 894 27303 900 27355
rect 1548 27303 1554 27355
rect 894 27183 1554 27303
rect 894 27131 900 27183
rect 1548 27131 1554 27183
rect 894 27011 1554 27131
rect 894 26959 900 27011
rect 1548 26959 1554 27011
rect 894 26839 1554 26959
rect 894 26787 900 26839
rect 1548 26787 1554 26839
rect 894 26667 1554 26787
rect 894 26615 900 26667
rect 1548 26615 1554 26667
rect 894 26495 1554 26615
rect 894 26443 900 26495
rect 1548 26443 1554 26495
rect 894 26323 1554 26443
rect 894 26271 900 26323
rect 1548 26271 1554 26323
rect 894 26151 1554 26271
rect 894 26099 900 26151
rect 1548 26099 1554 26151
rect 894 25979 1554 26099
rect 894 25927 900 25979
rect 1548 25927 1554 25979
rect 894 25807 1554 25927
rect 894 25755 900 25807
rect 1548 25755 1554 25807
rect 894 25635 1554 25755
rect 894 25583 900 25635
rect 1548 25583 1554 25635
rect 894 25463 1554 25583
rect 894 25411 900 25463
rect 1548 25411 1554 25463
rect 894 25291 1554 25411
rect 894 25239 900 25291
rect 1548 25239 1554 25291
rect 894 25119 1554 25239
rect 894 25067 900 25119
rect 1548 25067 1554 25119
rect 894 24947 1554 25067
rect 894 24895 900 24947
rect 1548 24895 1554 24947
rect 894 24775 1554 24895
rect 894 24723 900 24775
rect 1548 24723 1554 24775
rect 894 24603 1554 24723
rect 894 24551 900 24603
rect 1548 24551 1554 24603
rect 894 24431 1554 24551
rect 894 24379 900 24431
rect 1548 24379 1554 24431
rect 894 24259 1554 24379
rect 894 24207 900 24259
rect 1548 24207 1554 24259
rect 894 24087 1554 24207
rect 894 24035 900 24087
rect 1548 24035 1554 24087
rect 894 23915 1554 24035
rect 894 23863 900 23915
rect 1548 23863 1554 23915
rect 894 23743 1554 23863
rect 894 23691 900 23743
rect 1548 23691 1554 23743
rect 894 23571 1554 23691
rect 894 23519 900 23571
rect 1548 23519 1554 23571
rect 894 23399 1554 23519
rect 894 23347 900 23399
rect 1548 23347 1554 23399
rect 894 23227 1554 23347
rect 894 23175 900 23227
rect 1548 23175 1554 23227
rect 894 23055 1554 23175
rect 894 23003 900 23055
rect 1548 23003 1554 23055
rect 894 22883 1554 23003
rect 894 22831 900 22883
rect 1548 22831 1554 22883
rect 894 22711 1554 22831
rect 894 22659 900 22711
rect 1548 22659 1554 22711
rect 894 22539 1554 22659
rect 894 22487 900 22539
rect 1548 22487 1554 22539
rect 894 22367 1554 22487
rect 894 22315 900 22367
rect 1548 22315 1554 22367
rect 894 22195 1554 22315
rect 894 22143 900 22195
rect 1548 22143 1554 22195
rect 894 22023 1554 22143
rect 894 21971 900 22023
rect 1548 21971 1554 22023
rect 894 21851 1554 21971
rect 894 21799 900 21851
rect 1548 21799 1554 21851
rect 894 21679 1554 21799
rect 894 21627 900 21679
rect 1548 21627 1554 21679
rect 894 21507 1554 21627
rect 894 21455 900 21507
rect 1548 21455 1554 21507
rect 894 21335 1554 21455
rect 894 21283 900 21335
rect 1548 21283 1554 21335
rect 894 21163 1554 21283
rect 894 21111 900 21163
rect 1548 21111 1554 21163
rect 894 20991 1554 21111
rect 894 20939 900 20991
rect 1548 20939 1554 20991
rect 894 20819 1554 20939
rect 894 20767 900 20819
rect 1548 20767 1554 20819
rect 894 20647 1554 20767
rect 894 20595 900 20647
rect 1548 20595 1554 20647
rect 894 20475 1554 20595
rect 894 20423 900 20475
rect 1548 20423 1554 20475
rect 894 20303 1554 20423
rect 894 20251 900 20303
rect 1548 20251 1554 20303
rect 894 20131 1554 20251
rect 894 20079 900 20131
rect 1548 20079 1554 20131
rect 894 19959 1554 20079
rect 894 19907 900 19959
rect 1548 19907 1554 19959
rect 894 19787 1554 19907
rect 894 19735 900 19787
rect 1548 19735 1554 19787
rect 894 19615 1554 19735
rect 894 19563 900 19615
rect 1548 19563 1554 19615
rect 894 19443 1554 19563
rect 894 19391 900 19443
rect 1548 19391 1554 19443
rect 894 19271 1554 19391
rect 894 19219 900 19271
rect 1548 19219 1554 19271
rect 894 19099 1554 19219
rect 894 19047 900 19099
rect 1548 19047 1554 19099
rect 894 18927 1554 19047
rect 894 18875 900 18927
rect 1548 18875 1554 18927
rect 894 18755 1554 18875
rect 894 18703 900 18755
rect 1548 18703 1554 18755
rect 894 18583 1554 18703
rect 894 18531 900 18583
rect 1548 18531 1554 18583
rect 894 18411 1554 18531
rect 894 18359 900 18411
rect 1548 18359 1554 18411
rect 894 18239 1554 18359
rect 894 18187 900 18239
rect 1548 18187 1554 18239
rect 894 18067 1554 18187
rect 894 18015 900 18067
rect 1548 18015 1554 18067
rect 894 17895 1554 18015
rect 894 17843 900 17895
rect 1548 17843 1554 17895
rect 894 17723 1554 17843
rect 894 17671 900 17723
rect 1548 17671 1554 17723
rect 894 17551 1554 17671
rect 894 17499 900 17551
rect 1548 17499 1554 17551
rect 894 17379 1554 17499
rect 894 17327 900 17379
rect 1548 17327 1554 17379
rect 894 17207 1554 17327
rect 894 17155 900 17207
rect 1548 17155 1554 17207
rect 894 17035 1554 17155
rect 894 16983 900 17035
rect 1548 16983 1554 17035
rect 894 16863 1554 16983
rect 894 16811 900 16863
rect 1548 16811 1554 16863
rect 894 16691 1554 16811
rect 894 16639 900 16691
rect 1548 16639 1554 16691
rect 894 16519 1554 16639
rect 894 16467 900 16519
rect 1548 16467 1554 16519
rect 894 16347 1554 16467
rect 894 16295 900 16347
rect 1548 16295 1554 16347
rect 894 16175 1554 16295
rect 894 16123 900 16175
rect 1548 16123 1554 16175
rect 894 16003 1554 16123
rect 894 15951 900 16003
rect 1548 15951 1554 16003
rect 894 15831 1554 15951
rect 894 15779 900 15831
rect 1548 15779 1554 15831
rect 894 15659 1554 15779
rect 894 15607 900 15659
rect 1548 15607 1554 15659
rect 894 15487 1554 15607
rect 894 15435 900 15487
rect 1548 15435 1554 15487
rect 894 15315 1554 15435
rect 894 15263 900 15315
rect 1548 15263 1554 15315
rect 894 15143 1554 15263
rect 894 15091 900 15143
rect 1548 15091 1554 15143
rect 894 14971 1554 15091
rect 894 14919 900 14971
rect 1548 14919 1554 14971
rect 894 14799 1554 14919
rect 894 14747 900 14799
rect 1548 14747 1554 14799
rect 894 14627 1554 14747
rect 894 14575 900 14627
rect 1548 14575 1554 14627
rect 894 14455 1554 14575
rect 894 14403 900 14455
rect 1548 14403 1554 14455
rect 894 14283 1554 14403
rect 894 14231 900 14283
rect 1548 14231 1554 14283
rect 894 14111 1554 14231
rect 894 14059 900 14111
rect 1548 14059 1554 14111
rect 894 13939 1554 14059
rect 894 13887 900 13939
rect 1548 13887 1554 13939
rect 894 13767 1554 13887
rect 894 13715 900 13767
rect 1548 13715 1554 13767
rect 894 13595 1554 13715
rect 894 13543 900 13595
rect 1548 13543 1554 13595
rect 894 13423 1554 13543
rect 894 13371 900 13423
rect 1548 13371 1554 13423
rect 894 13251 1554 13371
rect 894 13199 900 13251
rect 1548 13199 1554 13251
rect 894 13079 1554 13199
rect 894 13027 900 13079
rect 1548 13027 1554 13079
rect 894 12907 1554 13027
rect 894 12855 900 12907
rect 1548 12855 1554 12907
rect 894 12735 1554 12855
rect 894 12683 900 12735
rect 1548 12683 1554 12735
rect 894 12563 1554 12683
rect 894 12511 900 12563
rect 1548 12511 1554 12563
rect 894 12391 1554 12511
rect 894 12339 900 12391
rect 1548 12339 1554 12391
rect 894 12219 1554 12339
rect 894 12167 900 12219
rect 1548 12167 1554 12219
rect 894 12047 1554 12167
rect 894 11995 900 12047
rect 1548 11995 1554 12047
rect 894 11875 1554 11995
rect 894 11823 900 11875
rect 1548 11823 1554 11875
rect 894 11703 1554 11823
rect 894 11651 900 11703
rect 1548 11651 1554 11703
rect 894 11531 1554 11651
rect 894 11479 900 11531
rect 1548 11479 1554 11531
rect 894 11359 1554 11479
rect 894 11307 900 11359
rect 1548 11307 1554 11359
rect 894 11187 1554 11307
rect 894 11135 900 11187
rect 1548 11135 1554 11187
rect 894 11015 1554 11135
rect 894 10963 900 11015
rect 1548 10963 1554 11015
rect 894 10843 1554 10963
rect 894 10791 900 10843
rect 1548 10791 1554 10843
rect 894 10671 1554 10791
rect 894 10619 900 10671
rect 1548 10619 1554 10671
rect 894 10499 1554 10619
rect 894 10447 900 10499
rect 1548 10447 1554 10499
rect 894 10327 1554 10447
rect 894 10275 900 10327
rect 1548 10275 1554 10327
rect 894 10155 1554 10275
rect 894 10103 900 10155
rect 1548 10103 1554 10155
rect 894 9983 1554 10103
rect 894 9931 900 9983
rect 1548 9931 1554 9983
rect 894 9811 1554 9931
rect 894 9759 900 9811
rect 1548 9759 1554 9811
rect 894 9639 1554 9759
rect 894 9587 900 9639
rect 1548 9587 1554 9639
rect 894 9467 1554 9587
rect 894 9415 900 9467
rect 1548 9415 1554 9467
rect 894 9295 1554 9415
rect 894 9243 900 9295
rect 1548 9243 1554 9295
rect 894 9123 1554 9243
rect 894 9071 900 9123
rect 1548 9071 1554 9123
rect 894 8951 1554 9071
rect 894 8899 900 8951
rect 1548 8899 1554 8951
rect 894 8779 1554 8899
rect 894 8727 900 8779
rect 1548 8727 1554 8779
rect 894 8607 1554 8727
rect 894 8555 900 8607
rect 1548 8555 1554 8607
rect 894 8435 1554 8555
rect 894 8383 900 8435
rect 1548 8383 1554 8435
rect 894 8263 1554 8383
rect 894 8211 900 8263
rect 1548 8211 1554 8263
rect 894 8091 1554 8211
rect 894 8039 900 8091
rect 1548 8039 1554 8091
rect 894 7919 1554 8039
rect 894 7867 900 7919
rect 1548 7867 1554 7919
rect 894 7747 1554 7867
rect 894 7695 900 7747
rect 1548 7695 1554 7747
rect 894 7575 1554 7695
rect 894 7523 900 7575
rect 1548 7523 1554 7575
rect 894 7403 1554 7523
rect 894 7351 900 7403
rect 1548 7351 1554 7403
rect 894 7231 1554 7351
rect 894 7179 900 7231
rect 1548 7179 1554 7231
rect 894 7059 1554 7179
rect 894 7007 900 7059
rect 1548 7007 1554 7059
rect 894 6887 1554 7007
rect 894 6835 900 6887
rect 1548 6835 1554 6887
rect 894 6715 1554 6835
rect 894 6663 900 6715
rect 1548 6663 1554 6715
rect 894 6543 1554 6663
rect 894 6491 900 6543
rect 1548 6491 1554 6543
rect 894 6371 1554 6491
rect 894 6319 900 6371
rect 1548 6319 1554 6371
rect 894 6199 1554 6319
rect 894 6147 900 6199
rect 1548 6147 1554 6199
rect 894 6027 1554 6147
rect 894 5975 900 6027
rect 1548 5975 1554 6027
rect 894 5855 1554 5975
rect 894 5803 900 5855
rect 1548 5803 1554 5855
rect 894 5683 1554 5803
rect 894 5631 900 5683
rect 1548 5631 1554 5683
rect 894 5511 1554 5631
rect 894 5459 900 5511
rect 1548 5459 1554 5511
rect 894 5339 1554 5459
rect 894 5287 900 5339
rect 1548 5287 1554 5339
rect 894 5167 1554 5287
rect 894 5115 900 5167
rect 1548 5115 1554 5167
rect 894 4995 1554 5115
rect 894 4943 900 4995
rect 1548 4943 1554 4995
rect 894 4823 1554 4943
rect 894 4771 900 4823
rect 1548 4771 1554 4823
rect 894 4651 1554 4771
rect 894 4599 900 4651
rect 1548 4599 1554 4651
rect 894 4479 1554 4599
rect 894 4427 900 4479
rect 1548 4427 1554 4479
rect 894 4307 1554 4427
rect 894 4255 900 4307
rect 1548 4255 1554 4307
rect 894 4135 1554 4255
rect 894 4083 900 4135
rect 1548 4083 1554 4135
rect 894 3963 1554 4083
rect 894 3911 900 3963
rect 1548 3911 1554 3963
rect 894 3791 1554 3911
rect 894 3739 900 3791
rect 1548 3739 1554 3791
rect 894 3619 1554 3739
rect 894 3567 900 3619
rect 1548 3567 1554 3619
rect 894 3447 1554 3567
rect 894 3395 900 3447
rect 1548 3395 1554 3447
rect 894 3275 1554 3395
rect 894 3223 900 3275
rect 1548 3223 1554 3275
rect 894 3103 1554 3223
rect 894 3051 900 3103
rect 1548 3051 1554 3103
rect 894 2931 1554 3051
rect 894 2879 900 2931
rect 1548 2879 1554 2931
rect 894 2759 1554 2879
rect 894 2707 900 2759
rect 1548 2707 1554 2759
rect 894 2587 1554 2707
rect 894 2535 900 2587
rect 1548 2535 1554 2587
rect 894 2415 1554 2535
rect 894 2363 900 2415
rect 1548 2363 1554 2415
rect 894 2243 1554 2363
rect 894 2191 900 2243
rect 1548 2191 1554 2243
rect 894 2071 1554 2191
rect 894 2019 900 2071
rect 1548 2019 1554 2071
rect 894 1899 1554 2019
rect 894 1847 900 1899
rect 1548 1847 1554 1899
rect 894 1727 1554 1847
rect 894 1675 900 1727
rect 1548 1675 1554 1727
rect 894 1555 1554 1675
rect 894 1503 900 1555
rect 1548 1503 1554 1555
rect 894 1383 1554 1503
rect 894 1331 900 1383
rect 1548 1331 1554 1383
rect 894 1211 1554 1331
rect 894 1159 900 1211
rect 1548 1159 1554 1211
rect 894 1039 1554 1159
rect 894 987 900 1039
rect 1548 987 1554 1039
rect 894 867 1554 987
rect 894 815 900 867
rect 1548 815 1554 867
rect 894 695 1554 815
rect 894 643 900 695
rect 1548 643 1554 695
rect 894 523 1554 643
rect 894 471 900 523
rect 1548 471 1554 523
rect 894 351 1554 471
rect 894 299 900 351
rect 1548 299 1554 351
rect 894 179 1554 299
rect 894 127 900 179
rect 1548 127 1554 179
rect 1618 43825 1672 43831
rect 1618 163 1672 169
<< end >>
