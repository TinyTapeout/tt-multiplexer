module vccd1_connection ();
endmodule