magic
tech sky130A
magscale 1 2
timestamp 1718271279
<< metal2 >>
rect 256 1115 916 1120
rect 256 5 265 1115
rect 907 5 916 1115
rect 256 0 916 5
rect 994 1115 1654 1120
rect 994 5 1089 1115
rect 1645 5 1654 1115
rect 994 0 1654 5
<< via2 >>
rect 265 5 907 1115
rect 1089 5 1645 1115
<< metal3 >>
rect 256 1119 960 1120
rect 256 1115 346 1119
rect 256 5 265 1115
rect 256 1 346 5
rect 954 1 960 1119
rect 256 0 960 1
rect 1080 1119 1840 1120
rect 1080 1115 1146 1119
rect 1080 5 1089 1115
rect 1080 1 1146 5
rect 1834 1 1840 1119
rect 1080 0 1840 1
<< via3 >>
rect 346 1115 954 1119
rect 346 5 907 1115
rect 907 5 954 1115
rect 346 1 954 5
rect 1146 1115 1834 1119
rect 1146 5 1645 1115
rect 1645 5 1834 1115
rect 1146 1 1834 5
<< metal4 >>
rect 0 0 240 1120
rect 340 1119 1040 1120
rect 340 1 346 1119
rect 954 1 1040 1119
rect 340 0 1040 1
rect 1140 1119 1840 1120
rect 1140 1 1146 1119
rect 1834 1 1840 1119
rect 1140 0 1840 1
<< end >>
