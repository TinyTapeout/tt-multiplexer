VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_pg_vdd_1
  CLASS BLOCK ;
  FOREIGN tt_pg_vdd_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.200 BY 111.520 ;
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000 0.000 1.200 110.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 8.000 0.000 9.200 110.000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.700 0.000 4.350 110.000 ;
    END
  END VPWR
  PIN GPWR
    DIRECTION OUTPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 4.850 0.000 7.500 110.000 ;
    END
  END GPWR
  PIN ctrl
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 231.000000 ;
    PORT
      LAYER met4 ;
        RECT 0.000 111.020 9.200 111.520 ;
    END
  END ctrl
  OBS
      LAYER nwell ;
        RECT 0.000 2.450 9.190 109.720 ;
      LAYER li1 ;
        RECT 0.180 2.630 9.010 109.660 ;
      LAYER met1 ;
        RECT 0.150 2.940 9.040 111.520 ;
      LAYER met2 ;
        RECT 0.150 3.070 9.040 111.480 ;
      LAYER met3 ;
        RECT 0.610 3.070 8.580 111.455 ;
  END
END tt_pg_vdd_1
END LIBRARY

