magic
tech sky130A
timestamp 1718083762
<< pwell >>
rect 6 0 914 212
<< nmos >>
rect 100 92 150 142
rect 190 92 240 142
rect 280 92 330 142
rect 370 92 420 142
rect 500 92 550 142
rect 590 92 640 142
rect 680 92 730 142
rect 770 92 820 142
<< ndiff >>
rect 63 151 92 155
rect 63 61 69 151
rect 86 142 92 151
rect 428 151 492 155
rect 428 142 434 151
rect 86 92 100 142
rect 150 92 190 142
rect 240 92 280 142
rect 330 92 370 142
rect 420 96 434 142
rect 486 142 492 151
rect 828 151 857 155
rect 828 142 834 151
rect 486 96 500 142
rect 420 92 500 96
rect 550 92 590 142
rect 640 92 680 142
rect 730 92 770 142
rect 820 92 834 142
rect 86 61 92 92
rect 63 57 92 61
rect 828 61 834 92
rect 851 61 857 151
rect 828 57 857 61
<< ndiffc >>
rect 69 61 86 151
rect 434 96 486 151
rect 834 61 851 151
<< psubdiff >>
rect 19 182 51 199
rect 869 182 901 199
rect 19 167 36 182
rect 884 167 901 182
rect 19 30 36 45
rect 884 30 901 45
rect 19 13 51 30
rect 869 13 901 30
<< psubdiffcont >>
rect 51 182 869 199
rect 19 45 36 167
rect 884 45 901 167
rect 51 13 869 30
<< poly >>
rect 100 142 150 155
rect 190 142 240 155
rect 280 142 330 155
rect 370 142 420 155
rect 500 142 550 155
rect 590 142 640 155
rect 680 142 730 155
rect 770 142 820 155
rect 100 76 150 92
rect 190 76 240 92
rect 280 76 330 92
rect 370 76 420 92
rect 500 76 550 92
rect 590 76 640 92
rect 680 76 730 92
rect 770 76 820 92
rect 100 71 820 76
rect 100 54 119 71
rect 803 54 820 71
rect 100 49 820 54
<< polycont >>
rect 119 54 803 71
<< locali >>
rect 19 182 51 199
rect 869 182 901 199
rect 19 167 36 182
rect 884 167 901 182
rect 428 156 492 159
rect 428 95 431 156
rect 489 95 492 156
rect 428 88 492 95
rect 111 54 119 71
rect 803 54 811 71
rect 19 30 36 45
rect 884 30 901 45
rect 19 13 51 30
rect 869 13 901 30
<< viali >>
rect 51 182 869 199
rect 19 45 36 167
rect 63 151 92 159
rect 63 61 69 151
rect 69 61 86 151
rect 86 61 92 151
rect 431 151 489 156
rect 431 96 434 151
rect 434 96 486 151
rect 486 96 489 151
rect 431 95 489 96
rect 828 151 857 159
rect 63 53 92 61
rect 119 54 803 71
rect 828 61 834 151
rect 834 61 851 151
rect 851 61 857 151
rect 828 53 857 61
rect 884 45 901 167
rect 51 13 869 30
<< metal1 >>
rect 16 199 904 202
rect 16 182 51 199
rect 869 182 904 199
rect 16 179 904 182
rect 16 167 95 179
rect 16 45 19 167
rect 36 159 95 167
rect 825 167 904 179
rect 36 53 63 159
rect 92 53 95 159
rect 425 102 428 161
rect 492 102 495 161
rect 425 95 431 102
rect 489 95 495 102
rect 425 92 495 95
rect 825 159 884 167
rect 36 45 95 53
rect 111 51 114 77
rect 367 74 370 77
rect 552 74 555 77
rect 367 71 555 74
rect 367 51 555 54
rect 808 51 811 77
rect 825 53 828 159
rect 857 53 884 159
rect 16 33 95 45
rect 825 45 884 53
rect 901 45 904 167
rect 825 33 904 45
rect 16 30 904 33
rect 16 13 51 30
rect 869 13 904 30
rect 16 10 904 13
<< via1 >>
rect 428 156 492 161
rect 428 102 431 156
rect 431 102 489 156
rect 489 102 492 156
rect 114 71 367 77
rect 555 71 808 77
rect 114 54 119 71
rect 119 54 367 71
rect 555 54 803 71
rect 803 54 808 71
rect 114 51 367 54
rect 555 51 808 54
<< metal2 >>
rect 425 102 428 161
rect 492 102 495 161
rect 111 51 114 77
rect 367 51 555 77
rect 808 51 811 77
<< properties >>
string FIXED_BBOX 0 0 920 212
<< end >>
