magic
tech sky130A
timestamp 1718199492
<< pwell >>
rect 6 0 914 262
<< nmos >>
rect 100 92 150 192
rect 190 92 240 192
rect 280 92 330 192
rect 370 92 420 192
rect 500 92 550 192
rect 590 92 640 192
rect 680 92 730 192
rect 770 92 820 192
<< ndiff >>
rect 63 201 92 205
rect 63 61 69 201
rect 86 192 92 201
rect 428 201 492 205
rect 428 192 434 201
rect 86 92 100 192
rect 150 92 190 192
rect 240 92 280 192
rect 330 92 370 192
rect 420 96 434 192
rect 486 192 492 201
rect 828 201 857 205
rect 828 192 834 201
rect 486 96 500 192
rect 420 92 500 96
rect 550 92 590 192
rect 640 92 680 192
rect 730 92 770 192
rect 820 92 834 192
rect 86 61 92 92
rect 63 57 92 61
rect 828 61 834 92
rect 851 61 857 201
rect 828 57 857 61
<< ndiffc >>
rect 69 61 86 201
rect 434 96 486 201
rect 834 61 851 201
<< psubdiff >>
rect 19 232 51 249
rect 869 232 901 249
rect 19 217 36 232
rect 884 217 901 232
rect 19 30 36 45
rect 884 30 901 45
rect 19 13 51 30
rect 869 13 901 30
<< psubdiffcont >>
rect 51 232 869 249
rect 19 45 36 217
rect 884 45 901 217
rect 51 13 869 30
<< poly >>
rect 100 192 150 205
rect 190 192 240 205
rect 280 192 330 205
rect 370 192 420 205
rect 500 192 550 205
rect 590 192 640 205
rect 680 192 730 205
rect 770 192 820 205
rect 100 76 150 92
rect 190 76 240 92
rect 280 76 330 92
rect 370 76 420 92
rect 500 76 550 92
rect 590 76 640 92
rect 680 76 730 92
rect 770 76 820 92
rect 100 71 820 76
rect 100 54 119 71
rect 803 54 820 71
rect 100 49 820 54
<< polycont >>
rect 119 54 803 71
<< locali >>
rect 19 232 51 249
rect 869 232 901 249
rect 19 217 36 232
rect 884 217 901 232
rect 428 206 492 209
rect 428 95 431 206
rect 489 95 492 206
rect 428 88 492 95
rect 111 54 119 71
rect 803 54 811 71
rect 19 30 36 45
rect 884 30 901 45
rect 19 13 51 30
rect 869 13 901 30
<< viali >>
rect 51 232 869 249
rect 19 45 36 217
rect 63 201 92 209
rect 63 61 69 201
rect 69 61 86 201
rect 86 61 92 201
rect 431 201 489 206
rect 431 96 434 201
rect 434 96 486 201
rect 486 96 489 201
rect 431 95 489 96
rect 828 201 857 209
rect 63 53 92 61
rect 119 54 803 71
rect 828 61 834 201
rect 834 61 851 201
rect 851 61 857 201
rect 828 53 857 61
rect 884 45 901 217
rect 51 13 869 30
<< metal1 >>
rect 16 249 904 252
rect 16 232 51 249
rect 869 232 904 249
rect 16 229 904 232
rect 16 217 95 229
rect 16 45 19 217
rect 36 209 95 217
rect 825 217 904 229
rect 36 53 63 209
rect 92 53 95 209
rect 425 102 428 211
rect 492 102 495 211
rect 425 95 431 102
rect 489 95 495 102
rect 425 92 495 95
rect 825 209 884 217
rect 36 45 95 53
rect 111 51 114 77
rect 367 74 370 77
rect 552 74 555 77
rect 367 71 555 74
rect 367 51 555 54
rect 808 51 811 77
rect 825 53 828 209
rect 857 53 884 209
rect 16 33 95 45
rect 825 45 884 53
rect 901 45 904 217
rect 825 33 904 45
rect 16 30 904 33
rect 16 13 51 30
rect 869 13 904 30
rect 16 10 904 13
<< via1 >>
rect 428 206 492 211
rect 428 102 431 206
rect 431 102 489 206
rect 489 102 492 206
rect 114 71 367 77
rect 555 71 808 77
rect 114 54 119 71
rect 119 54 367 71
rect 555 54 803 71
rect 803 54 808 71
rect 114 51 367 54
rect 555 51 808 54
<< metal2 >>
rect 425 102 428 211
rect 492 102 495 211
rect 111 51 114 77
rect 367 51 555 77
rect 808 51 811 77
<< properties >>
string FIXED_BBOX 0 0 920 262
<< end >>
