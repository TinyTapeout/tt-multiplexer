** sch_path: /home/tnt/consult/tinytapeout/tt-multiplexer/pg/tt_pg_1v8_2/xschem/tt_pg_1v8_2.sch
.subckt tt_pg_1v8_2 VGND VPWR ctrl GPWR
*.PININFO ctrl:I VGND:B VPWR:B GPWR:B
XM2 ctrl_n ctrl VGND VGND sky130_fd_pr__nfet_01v8 L=0.15 W=3.5 nf=2 m=1
XM1 ctrl_n ctrl VPWR VPWR sky130_fd_pr__pfet_01v8_hvt L=0.15 W=10.5 nf=2 m=1
XM3 GPWR ctrl_n VPWR VPWR sky130_fd_pr__pfet_01v8 L=0.15 W=3683 nf=508 m=1
XM4 GPWR ctrl_n net1 VGND sky130_fd_pr__nfet_01v8 L=0.5 W=1 nf=1 m=1
XM5 net1 ctrl_n net2 VGND sky130_fd_pr__nfet_01v8 L=0.5 W=1 nf=1 m=1
XM6 net2 ctrl_n net3 VGND sky130_fd_pr__nfet_01v8 L=0.5 W=1 nf=1 m=1
XM7 net3 ctrl_n VGND VGND sky130_fd_pr__nfet_01v8 L=0.5 W=1 nf=1 m=1
XM8 GPWR ctrl_n net4 VGND sky130_fd_pr__nfet_01v8 L=0.5 W=1 nf=1 m=1
XM9 net4 ctrl_n net5 VGND sky130_fd_pr__nfet_01v8 L=0.5 W=1 nf=1 m=1
XM10 net5 ctrl_n net6 VGND sky130_fd_pr__nfet_01v8 L=0.5 W=1 nf=1 m=1
XM11 net6 ctrl_n VGND VGND sky130_fd_pr__nfet_01v8 L=0.5 W=1 nf=1 m=1
XC1 VPWR VGND sky130_fd_pr__cap_mim_m3_1 W=6.9 L=19.4 m=2
XC2 GPWR VGND sky130_fd_pr__cap_mim_m3_1 W=6.9 L=19.4 m=4
.ends
.end
