magic
tech sky130A
timestamp 1710930057
<< checkpaint >>
rect -570 546 2410 2806
rect -570 -630 810 546
rect 1030 -630 2410 546
<< metal3 >>
rect 60 2173 180 2176
rect 60 1179 63 2173
rect 177 1179 180 2173
rect 445 2086 475 2176
rect 875 2173 965 2176
rect 875 1979 878 2173
rect 962 1979 965 2173
rect 875 1976 965 1979
rect 1660 2173 1780 2176
rect 60 1176 180 1179
rect 875 1373 965 1376
rect 875 1179 878 1373
rect 962 1179 965 1373
rect 875 1176 965 1179
rect 1660 1179 1663 2173
rect 1777 1179 1780 2173
rect 1660 1176 1780 1179
<< via3 >>
rect 63 1179 177 2173
rect 878 1979 962 2173
rect 878 1179 962 1373
rect 1663 1179 1777 2173
<< metal4 >>
rect 60 2173 180 2176
rect 60 1179 63 2173
rect 177 1179 180 2173
rect 875 2173 965 2176
rect 875 1979 878 2173
rect 962 1979 965 2173
rect 875 1976 965 1979
rect 1660 2173 1780 2176
rect 60 0 180 1179
rect 875 1373 965 1376
rect 875 1179 878 1373
rect 962 1179 965 1373
rect 875 1176 965 1179
rect 1660 1179 1663 2173
rect 1777 1179 1780 2173
rect 1660 0 1780 1179
<< labels >>
rlabel metal4 60 0 180 2176 1 VGND
port 1 n ground input
rlabel metal4 1660 0 1780 2176 1 VPWR
port 2 n power input
rlabel metal4 875 1976 965 2176 1 mod
port 3 n analog bidirectional
rlabel metal4 875 1176 965 1376 1 bus
port 4 n analog bidirectional
rlabel metal3 445 2086 475 2176 1 ctrl
port 5 n signal input
<< properties >>
string FIXED_BBOX 0 0 1840 2176
<< end >>
