magic
tech sky130A
magscale 1 2
timestamp 1697797911
<< nwell >>
rect 0 22898 1838 44352
rect 0 400 1838 21854
<< pmos >>
rect 219 44122 1619 44152
rect 219 44026 1619 44056
rect 219 43930 1619 43960
rect 219 43834 1619 43864
rect 219 43738 1619 43768
rect 219 43642 1619 43672
rect 219 43546 1619 43576
rect 219 43450 1619 43480
rect 219 43354 1619 43384
rect 219 43258 1619 43288
rect 219 43162 1619 43192
rect 219 43066 1619 43096
rect 219 42970 1619 43000
rect 219 42874 1619 42904
rect 219 42778 1619 42808
rect 219 42682 1619 42712
rect 219 42586 1619 42616
rect 219 42490 1619 42520
rect 219 42394 1619 42424
rect 219 42298 1619 42328
rect 219 42202 1619 42232
rect 219 42106 1619 42136
rect 219 42010 1619 42040
rect 219 41914 1619 41944
rect 219 41818 1619 41848
rect 219 41722 1619 41752
rect 219 41626 1619 41656
rect 219 41530 1619 41560
rect 219 41434 1619 41464
rect 219 41338 1619 41368
rect 219 41242 1619 41272
rect 219 41146 1619 41176
rect 219 41050 1619 41080
rect 219 40954 1619 40984
rect 219 40858 1619 40888
rect 219 40762 1619 40792
rect 219 40666 1619 40696
rect 219 40570 1619 40600
rect 219 40474 1619 40504
rect 219 40378 1619 40408
rect 219 40282 1619 40312
rect 219 40186 1619 40216
rect 219 40090 1619 40120
rect 219 39994 1619 40024
rect 219 39898 1619 39928
rect 219 39802 1619 39832
rect 219 39706 1619 39736
rect 219 39610 1619 39640
rect 219 39514 1619 39544
rect 219 39418 1619 39448
rect 219 39322 1619 39352
rect 219 39226 1619 39256
rect 219 39130 1619 39160
rect 219 39034 1619 39064
rect 219 38938 1619 38968
rect 219 38842 1619 38872
rect 219 38746 1619 38776
rect 219 38650 1619 38680
rect 219 38554 1619 38584
rect 219 38458 1619 38488
rect 219 38362 1619 38392
rect 219 38266 1619 38296
rect 219 38170 1619 38200
rect 219 38074 1619 38104
rect 219 37978 1619 38008
rect 219 37882 1619 37912
rect 219 37786 1619 37816
rect 219 37690 1619 37720
rect 219 37594 1619 37624
rect 219 37498 1619 37528
rect 219 37402 1619 37432
rect 219 37306 1619 37336
rect 219 37210 1619 37240
rect 219 37114 1619 37144
rect 219 37018 1619 37048
rect 219 36922 1619 36952
rect 219 36826 1619 36856
rect 219 36730 1619 36760
rect 219 36634 1619 36664
rect 219 36538 1619 36568
rect 219 36442 1619 36472
rect 219 36346 1619 36376
rect 219 36250 1619 36280
rect 219 36154 1619 36184
rect 219 36058 1619 36088
rect 219 35962 1619 35992
rect 219 35866 1619 35896
rect 219 35770 1619 35800
rect 219 35674 1619 35704
rect 219 35578 1619 35608
rect 219 35482 1619 35512
rect 219 35386 1619 35416
rect 219 35290 1619 35320
rect 219 35194 1619 35224
rect 219 35098 1619 35128
rect 219 35002 1619 35032
rect 219 34906 1619 34936
rect 219 34810 1619 34840
rect 219 34714 1619 34744
rect 219 34618 1619 34648
rect 219 34522 1619 34552
rect 219 34426 1619 34456
rect 219 34330 1619 34360
rect 219 34234 1619 34264
rect 219 34138 1619 34168
rect 219 34042 1619 34072
rect 219 33946 1619 33976
rect 219 33850 1619 33880
rect 219 33754 1619 33784
rect 219 33658 1619 33688
rect 219 33562 1619 33592
rect 219 33466 1619 33496
rect 219 33370 1619 33400
rect 219 33274 1619 33304
rect 219 33178 1619 33208
rect 219 33082 1619 33112
rect 219 32986 1619 33016
rect 219 32890 1619 32920
rect 219 32794 1619 32824
rect 219 32698 1619 32728
rect 219 32602 1619 32632
rect 219 32506 1619 32536
rect 219 32410 1619 32440
rect 219 32314 1619 32344
rect 219 32218 1619 32248
rect 219 32122 1619 32152
rect 219 32026 1619 32056
rect 219 31930 1619 31960
rect 219 31834 1619 31864
rect 219 31738 1619 31768
rect 219 31642 1619 31672
rect 219 31546 1619 31576
rect 219 31450 1619 31480
rect 219 31354 1619 31384
rect 219 31258 1619 31288
rect 219 31162 1619 31192
rect 219 31066 1619 31096
rect 219 30970 1619 31000
rect 219 30874 1619 30904
rect 219 30778 1619 30808
rect 219 30682 1619 30712
rect 219 30586 1619 30616
rect 219 30490 1619 30520
rect 219 30394 1619 30424
rect 219 30298 1619 30328
rect 219 30202 1619 30232
rect 219 30106 1619 30136
rect 219 30010 1619 30040
rect 219 29914 1619 29944
rect 219 29818 1619 29848
rect 219 29722 1619 29752
rect 219 29626 1619 29656
rect 219 29530 1619 29560
rect 219 29434 1619 29464
rect 219 29338 1619 29368
rect 219 29242 1619 29272
rect 219 29146 1619 29176
rect 219 29050 1619 29080
rect 219 28954 1619 28984
rect 219 28858 1619 28888
rect 219 28762 1619 28792
rect 219 28666 1619 28696
rect 219 28570 1619 28600
rect 219 28474 1619 28504
rect 219 28378 1619 28408
rect 219 28282 1619 28312
rect 219 28186 1619 28216
rect 219 28090 1619 28120
rect 219 27994 1619 28024
rect 219 27898 1619 27928
rect 219 27802 1619 27832
rect 219 27706 1619 27736
rect 219 27610 1619 27640
rect 219 27514 1619 27544
rect 219 27418 1619 27448
rect 219 27322 1619 27352
rect 219 27226 1619 27256
rect 219 27130 1619 27160
rect 219 27034 1619 27064
rect 219 26938 1619 26968
rect 219 26842 1619 26872
rect 219 26746 1619 26776
rect 219 26650 1619 26680
rect 219 26554 1619 26584
rect 219 26458 1619 26488
rect 219 26362 1619 26392
rect 219 26266 1619 26296
rect 219 26170 1619 26200
rect 219 26074 1619 26104
rect 219 25978 1619 26008
rect 219 25882 1619 25912
rect 219 25786 1619 25816
rect 219 25690 1619 25720
rect 219 25594 1619 25624
rect 219 25498 1619 25528
rect 219 25402 1619 25432
rect 219 25306 1619 25336
rect 219 25210 1619 25240
rect 219 25114 1619 25144
rect 219 25018 1619 25048
rect 219 24922 1619 24952
rect 219 24826 1619 24856
rect 219 24730 1619 24760
rect 219 24634 1619 24664
rect 219 24538 1619 24568
rect 219 24442 1619 24472
rect 219 24346 1619 24376
rect 219 24250 1619 24280
rect 219 24154 1619 24184
rect 219 24058 1619 24088
rect 219 23962 1619 23992
rect 219 23866 1619 23896
rect 219 23770 1619 23800
rect 219 23674 1619 23704
rect 219 23578 1619 23608
rect 219 23482 1619 23512
rect 219 23386 1619 23416
rect 219 23290 1619 23320
rect 219 23194 1619 23224
rect 219 23098 1619 23128
rect 219 21624 1619 21654
rect 219 21528 1619 21558
rect 219 21432 1619 21462
rect 219 21336 1619 21366
rect 219 21240 1619 21270
rect 219 21144 1619 21174
rect 219 21048 1619 21078
rect 219 20952 1619 20982
rect 219 20856 1619 20886
rect 219 20760 1619 20790
rect 219 20664 1619 20694
rect 219 20568 1619 20598
rect 219 20472 1619 20502
rect 219 20376 1619 20406
rect 219 20280 1619 20310
rect 219 20184 1619 20214
rect 219 20088 1619 20118
rect 219 19992 1619 20022
rect 219 19896 1619 19926
rect 219 19800 1619 19830
rect 219 19704 1619 19734
rect 219 19608 1619 19638
rect 219 19512 1619 19542
rect 219 19416 1619 19446
rect 219 19320 1619 19350
rect 219 19224 1619 19254
rect 219 19128 1619 19158
rect 219 19032 1619 19062
rect 219 18936 1619 18966
rect 219 18840 1619 18870
rect 219 18744 1619 18774
rect 219 18648 1619 18678
rect 219 18552 1619 18582
rect 219 18456 1619 18486
rect 219 18360 1619 18390
rect 219 18264 1619 18294
rect 219 18168 1619 18198
rect 219 18072 1619 18102
rect 219 17976 1619 18006
rect 219 17880 1619 17910
rect 219 17784 1619 17814
rect 219 17688 1619 17718
rect 219 17592 1619 17622
rect 219 17496 1619 17526
rect 219 17400 1619 17430
rect 219 17304 1619 17334
rect 219 17208 1619 17238
rect 219 17112 1619 17142
rect 219 17016 1619 17046
rect 219 16920 1619 16950
rect 219 16824 1619 16854
rect 219 16728 1619 16758
rect 219 16632 1619 16662
rect 219 16536 1619 16566
rect 219 16440 1619 16470
rect 219 16344 1619 16374
rect 219 16248 1619 16278
rect 219 16152 1619 16182
rect 219 16056 1619 16086
rect 219 15960 1619 15990
rect 219 15864 1619 15894
rect 219 15768 1619 15798
rect 219 15672 1619 15702
rect 219 15576 1619 15606
rect 219 15480 1619 15510
rect 219 15384 1619 15414
rect 219 15288 1619 15318
rect 219 15192 1619 15222
rect 219 15096 1619 15126
rect 219 15000 1619 15030
rect 219 14904 1619 14934
rect 219 14808 1619 14838
rect 219 14712 1619 14742
rect 219 14616 1619 14646
rect 219 14520 1619 14550
rect 219 14424 1619 14454
rect 219 14328 1619 14358
rect 219 14232 1619 14262
rect 219 14136 1619 14166
rect 219 14040 1619 14070
rect 219 13944 1619 13974
rect 219 13848 1619 13878
rect 219 13752 1619 13782
rect 219 13656 1619 13686
rect 219 13560 1619 13590
rect 219 13464 1619 13494
rect 219 13368 1619 13398
rect 219 13272 1619 13302
rect 219 13176 1619 13206
rect 219 13080 1619 13110
rect 219 12984 1619 13014
rect 219 12888 1619 12918
rect 219 12792 1619 12822
rect 219 12696 1619 12726
rect 219 12600 1619 12630
rect 219 12504 1619 12534
rect 219 12408 1619 12438
rect 219 12312 1619 12342
rect 219 12216 1619 12246
rect 219 12120 1619 12150
rect 219 12024 1619 12054
rect 219 11928 1619 11958
rect 219 11832 1619 11862
rect 219 11736 1619 11766
rect 219 11640 1619 11670
rect 219 11544 1619 11574
rect 219 11448 1619 11478
rect 219 11352 1619 11382
rect 219 11256 1619 11286
rect 219 11160 1619 11190
rect 219 11064 1619 11094
rect 219 10968 1619 10998
rect 219 10872 1619 10902
rect 219 10776 1619 10806
rect 219 10680 1619 10710
rect 219 10584 1619 10614
rect 219 10488 1619 10518
rect 219 10392 1619 10422
rect 219 10296 1619 10326
rect 219 10200 1619 10230
rect 219 10104 1619 10134
rect 219 10008 1619 10038
rect 219 9912 1619 9942
rect 219 9816 1619 9846
rect 219 9720 1619 9750
rect 219 9624 1619 9654
rect 219 9528 1619 9558
rect 219 9432 1619 9462
rect 219 9336 1619 9366
rect 219 9240 1619 9270
rect 219 9144 1619 9174
rect 219 9048 1619 9078
rect 219 8952 1619 8982
rect 219 8856 1619 8886
rect 219 8760 1619 8790
rect 219 8664 1619 8694
rect 219 8568 1619 8598
rect 219 8472 1619 8502
rect 219 8376 1619 8406
rect 219 8280 1619 8310
rect 219 8184 1619 8214
rect 219 8088 1619 8118
rect 219 7992 1619 8022
rect 219 7896 1619 7926
rect 219 7800 1619 7830
rect 219 7704 1619 7734
rect 219 7608 1619 7638
rect 219 7512 1619 7542
rect 219 7416 1619 7446
rect 219 7320 1619 7350
rect 219 7224 1619 7254
rect 219 7128 1619 7158
rect 219 7032 1619 7062
rect 219 6936 1619 6966
rect 219 6840 1619 6870
rect 219 6744 1619 6774
rect 219 6648 1619 6678
rect 219 6552 1619 6582
rect 219 6456 1619 6486
rect 219 6360 1619 6390
rect 219 6264 1619 6294
rect 219 6168 1619 6198
rect 219 6072 1619 6102
rect 219 5976 1619 6006
rect 219 5880 1619 5910
rect 219 5784 1619 5814
rect 219 5688 1619 5718
rect 219 5592 1619 5622
rect 219 5496 1619 5526
rect 219 5400 1619 5430
rect 219 5304 1619 5334
rect 219 5208 1619 5238
rect 219 5112 1619 5142
rect 219 5016 1619 5046
rect 219 4920 1619 4950
rect 219 4824 1619 4854
rect 219 4728 1619 4758
rect 219 4632 1619 4662
rect 219 4536 1619 4566
rect 219 4440 1619 4470
rect 219 4344 1619 4374
rect 219 4248 1619 4278
rect 219 4152 1619 4182
rect 219 4056 1619 4086
rect 219 3960 1619 3990
rect 219 3864 1619 3894
rect 219 3768 1619 3798
rect 219 3672 1619 3702
rect 219 3576 1619 3606
rect 219 3480 1619 3510
rect 219 3384 1619 3414
rect 219 3288 1619 3318
rect 219 3192 1619 3222
rect 219 3096 1619 3126
rect 219 3000 1619 3030
rect 219 2904 1619 2934
rect 219 2808 1619 2838
rect 219 2712 1619 2742
rect 219 2616 1619 2646
rect 219 2520 1619 2550
rect 219 2424 1619 2454
rect 219 2328 1619 2358
rect 219 2232 1619 2262
rect 219 2136 1619 2166
rect 219 2040 1619 2070
rect 219 1944 1619 1974
rect 219 1848 1619 1878
rect 219 1752 1619 1782
rect 219 1656 1619 1686
rect 219 1560 1619 1590
rect 219 1464 1619 1494
rect 219 1368 1619 1398
rect 219 1272 1619 1302
rect 219 1176 1619 1206
rect 219 1080 1619 1110
rect 219 984 1619 1014
rect 219 888 1619 918
rect 219 792 1619 822
rect 219 696 1619 726
rect 219 600 1619 630
<< pdiff >>
rect 219 44202 1619 44214
rect 219 44168 231 44202
rect 1607 44168 1619 44202
rect 219 44152 1619 44168
rect 219 44106 1619 44122
rect 219 44072 231 44106
rect 1607 44072 1619 44106
rect 219 44056 1619 44072
rect 219 44010 1619 44026
rect 219 43976 231 44010
rect 1607 43976 1619 44010
rect 219 43960 1619 43976
rect 219 43914 1619 43930
rect 219 43880 231 43914
rect 1607 43880 1619 43914
rect 219 43864 1619 43880
rect 219 43818 1619 43834
rect 219 43784 231 43818
rect 1607 43784 1619 43818
rect 219 43768 1619 43784
rect 219 43722 1619 43738
rect 219 43688 231 43722
rect 1607 43688 1619 43722
rect 219 43672 1619 43688
rect 219 43626 1619 43642
rect 219 43592 231 43626
rect 1607 43592 1619 43626
rect 219 43576 1619 43592
rect 219 43530 1619 43546
rect 219 43496 231 43530
rect 1607 43496 1619 43530
rect 219 43480 1619 43496
rect 219 43434 1619 43450
rect 219 43400 231 43434
rect 1607 43400 1619 43434
rect 219 43384 1619 43400
rect 219 43338 1619 43354
rect 219 43304 231 43338
rect 1607 43304 1619 43338
rect 219 43288 1619 43304
rect 219 43242 1619 43258
rect 219 43208 231 43242
rect 1607 43208 1619 43242
rect 219 43192 1619 43208
rect 219 43146 1619 43162
rect 219 43112 231 43146
rect 1607 43112 1619 43146
rect 219 43096 1619 43112
rect 219 43050 1619 43066
rect 219 43016 231 43050
rect 1607 43016 1619 43050
rect 219 43000 1619 43016
rect 219 42954 1619 42970
rect 219 42920 231 42954
rect 1607 42920 1619 42954
rect 219 42904 1619 42920
rect 219 42858 1619 42874
rect 219 42824 231 42858
rect 1607 42824 1619 42858
rect 219 42808 1619 42824
rect 219 42762 1619 42778
rect 219 42728 231 42762
rect 1607 42728 1619 42762
rect 219 42712 1619 42728
rect 219 42666 1619 42682
rect 219 42632 231 42666
rect 1607 42632 1619 42666
rect 219 42616 1619 42632
rect 219 42570 1619 42586
rect 219 42536 231 42570
rect 1607 42536 1619 42570
rect 219 42520 1619 42536
rect 219 42474 1619 42490
rect 219 42440 231 42474
rect 1607 42440 1619 42474
rect 219 42424 1619 42440
rect 219 42378 1619 42394
rect 219 42344 231 42378
rect 1607 42344 1619 42378
rect 219 42328 1619 42344
rect 219 42282 1619 42298
rect 219 42248 231 42282
rect 1607 42248 1619 42282
rect 219 42232 1619 42248
rect 219 42186 1619 42202
rect 219 42152 231 42186
rect 1607 42152 1619 42186
rect 219 42136 1619 42152
rect 219 42090 1619 42106
rect 219 42056 231 42090
rect 1607 42056 1619 42090
rect 219 42040 1619 42056
rect 219 41994 1619 42010
rect 219 41960 231 41994
rect 1607 41960 1619 41994
rect 219 41944 1619 41960
rect 219 41898 1619 41914
rect 219 41864 231 41898
rect 1607 41864 1619 41898
rect 219 41848 1619 41864
rect 219 41802 1619 41818
rect 219 41768 231 41802
rect 1607 41768 1619 41802
rect 219 41752 1619 41768
rect 219 41706 1619 41722
rect 219 41672 231 41706
rect 1607 41672 1619 41706
rect 219 41656 1619 41672
rect 219 41610 1619 41626
rect 219 41576 231 41610
rect 1607 41576 1619 41610
rect 219 41560 1619 41576
rect 219 41514 1619 41530
rect 219 41480 231 41514
rect 1607 41480 1619 41514
rect 219 41464 1619 41480
rect 219 41418 1619 41434
rect 219 41384 231 41418
rect 1607 41384 1619 41418
rect 219 41368 1619 41384
rect 219 41322 1619 41338
rect 219 41288 231 41322
rect 1607 41288 1619 41322
rect 219 41272 1619 41288
rect 219 41226 1619 41242
rect 219 41192 231 41226
rect 1607 41192 1619 41226
rect 219 41176 1619 41192
rect 219 41130 1619 41146
rect 219 41096 231 41130
rect 1607 41096 1619 41130
rect 219 41080 1619 41096
rect 219 41034 1619 41050
rect 219 41000 231 41034
rect 1607 41000 1619 41034
rect 219 40984 1619 41000
rect 219 40938 1619 40954
rect 219 40904 231 40938
rect 1607 40904 1619 40938
rect 219 40888 1619 40904
rect 219 40842 1619 40858
rect 219 40808 231 40842
rect 1607 40808 1619 40842
rect 219 40792 1619 40808
rect 219 40746 1619 40762
rect 219 40712 231 40746
rect 1607 40712 1619 40746
rect 219 40696 1619 40712
rect 219 40650 1619 40666
rect 219 40616 231 40650
rect 1607 40616 1619 40650
rect 219 40600 1619 40616
rect 219 40554 1619 40570
rect 219 40520 231 40554
rect 1607 40520 1619 40554
rect 219 40504 1619 40520
rect 219 40458 1619 40474
rect 219 40424 231 40458
rect 1607 40424 1619 40458
rect 219 40408 1619 40424
rect 219 40362 1619 40378
rect 219 40328 231 40362
rect 1607 40328 1619 40362
rect 219 40312 1619 40328
rect 219 40266 1619 40282
rect 219 40232 231 40266
rect 1607 40232 1619 40266
rect 219 40216 1619 40232
rect 219 40170 1619 40186
rect 219 40136 231 40170
rect 1607 40136 1619 40170
rect 219 40120 1619 40136
rect 219 40074 1619 40090
rect 219 40040 231 40074
rect 1607 40040 1619 40074
rect 219 40024 1619 40040
rect 219 39978 1619 39994
rect 219 39944 231 39978
rect 1607 39944 1619 39978
rect 219 39928 1619 39944
rect 219 39882 1619 39898
rect 219 39848 231 39882
rect 1607 39848 1619 39882
rect 219 39832 1619 39848
rect 219 39786 1619 39802
rect 219 39752 231 39786
rect 1607 39752 1619 39786
rect 219 39736 1619 39752
rect 219 39690 1619 39706
rect 219 39656 231 39690
rect 1607 39656 1619 39690
rect 219 39640 1619 39656
rect 219 39594 1619 39610
rect 219 39560 231 39594
rect 1607 39560 1619 39594
rect 219 39544 1619 39560
rect 219 39498 1619 39514
rect 219 39464 231 39498
rect 1607 39464 1619 39498
rect 219 39448 1619 39464
rect 219 39402 1619 39418
rect 219 39368 231 39402
rect 1607 39368 1619 39402
rect 219 39352 1619 39368
rect 219 39306 1619 39322
rect 219 39272 231 39306
rect 1607 39272 1619 39306
rect 219 39256 1619 39272
rect 219 39210 1619 39226
rect 219 39176 231 39210
rect 1607 39176 1619 39210
rect 219 39160 1619 39176
rect 219 39114 1619 39130
rect 219 39080 231 39114
rect 1607 39080 1619 39114
rect 219 39064 1619 39080
rect 219 39018 1619 39034
rect 219 38984 231 39018
rect 1607 38984 1619 39018
rect 219 38968 1619 38984
rect 219 38922 1619 38938
rect 219 38888 231 38922
rect 1607 38888 1619 38922
rect 219 38872 1619 38888
rect 219 38826 1619 38842
rect 219 38792 231 38826
rect 1607 38792 1619 38826
rect 219 38776 1619 38792
rect 219 38730 1619 38746
rect 219 38696 231 38730
rect 1607 38696 1619 38730
rect 219 38680 1619 38696
rect 219 38634 1619 38650
rect 219 38600 231 38634
rect 1607 38600 1619 38634
rect 219 38584 1619 38600
rect 219 38538 1619 38554
rect 219 38504 231 38538
rect 1607 38504 1619 38538
rect 219 38488 1619 38504
rect 219 38442 1619 38458
rect 219 38408 231 38442
rect 1607 38408 1619 38442
rect 219 38392 1619 38408
rect 219 38346 1619 38362
rect 219 38312 231 38346
rect 1607 38312 1619 38346
rect 219 38296 1619 38312
rect 219 38250 1619 38266
rect 219 38216 231 38250
rect 1607 38216 1619 38250
rect 219 38200 1619 38216
rect 219 38154 1619 38170
rect 219 38120 231 38154
rect 1607 38120 1619 38154
rect 219 38104 1619 38120
rect 219 38058 1619 38074
rect 219 38024 231 38058
rect 1607 38024 1619 38058
rect 219 38008 1619 38024
rect 219 37962 1619 37978
rect 219 37928 231 37962
rect 1607 37928 1619 37962
rect 219 37912 1619 37928
rect 219 37866 1619 37882
rect 219 37832 231 37866
rect 1607 37832 1619 37866
rect 219 37816 1619 37832
rect 219 37770 1619 37786
rect 219 37736 231 37770
rect 1607 37736 1619 37770
rect 219 37720 1619 37736
rect 219 37674 1619 37690
rect 219 37640 231 37674
rect 1607 37640 1619 37674
rect 219 37624 1619 37640
rect 219 37578 1619 37594
rect 219 37544 231 37578
rect 1607 37544 1619 37578
rect 219 37528 1619 37544
rect 219 37482 1619 37498
rect 219 37448 231 37482
rect 1607 37448 1619 37482
rect 219 37432 1619 37448
rect 219 37386 1619 37402
rect 219 37352 231 37386
rect 1607 37352 1619 37386
rect 219 37336 1619 37352
rect 219 37290 1619 37306
rect 219 37256 231 37290
rect 1607 37256 1619 37290
rect 219 37240 1619 37256
rect 219 37194 1619 37210
rect 219 37160 231 37194
rect 1607 37160 1619 37194
rect 219 37144 1619 37160
rect 219 37098 1619 37114
rect 219 37064 231 37098
rect 1607 37064 1619 37098
rect 219 37048 1619 37064
rect 219 37002 1619 37018
rect 219 36968 231 37002
rect 1607 36968 1619 37002
rect 219 36952 1619 36968
rect 219 36906 1619 36922
rect 219 36872 231 36906
rect 1607 36872 1619 36906
rect 219 36856 1619 36872
rect 219 36810 1619 36826
rect 219 36776 231 36810
rect 1607 36776 1619 36810
rect 219 36760 1619 36776
rect 219 36714 1619 36730
rect 219 36680 231 36714
rect 1607 36680 1619 36714
rect 219 36664 1619 36680
rect 219 36618 1619 36634
rect 219 36584 231 36618
rect 1607 36584 1619 36618
rect 219 36568 1619 36584
rect 219 36522 1619 36538
rect 219 36488 231 36522
rect 1607 36488 1619 36522
rect 219 36472 1619 36488
rect 219 36426 1619 36442
rect 219 36392 231 36426
rect 1607 36392 1619 36426
rect 219 36376 1619 36392
rect 219 36330 1619 36346
rect 219 36296 231 36330
rect 1607 36296 1619 36330
rect 219 36280 1619 36296
rect 219 36234 1619 36250
rect 219 36200 231 36234
rect 1607 36200 1619 36234
rect 219 36184 1619 36200
rect 219 36138 1619 36154
rect 219 36104 231 36138
rect 1607 36104 1619 36138
rect 219 36088 1619 36104
rect 219 36042 1619 36058
rect 219 36008 231 36042
rect 1607 36008 1619 36042
rect 219 35992 1619 36008
rect 219 35946 1619 35962
rect 219 35912 231 35946
rect 1607 35912 1619 35946
rect 219 35896 1619 35912
rect 219 35850 1619 35866
rect 219 35816 231 35850
rect 1607 35816 1619 35850
rect 219 35800 1619 35816
rect 219 35754 1619 35770
rect 219 35720 231 35754
rect 1607 35720 1619 35754
rect 219 35704 1619 35720
rect 219 35658 1619 35674
rect 219 35624 231 35658
rect 1607 35624 1619 35658
rect 219 35608 1619 35624
rect 219 35562 1619 35578
rect 219 35528 231 35562
rect 1607 35528 1619 35562
rect 219 35512 1619 35528
rect 219 35466 1619 35482
rect 219 35432 231 35466
rect 1607 35432 1619 35466
rect 219 35416 1619 35432
rect 219 35370 1619 35386
rect 219 35336 231 35370
rect 1607 35336 1619 35370
rect 219 35320 1619 35336
rect 219 35274 1619 35290
rect 219 35240 231 35274
rect 1607 35240 1619 35274
rect 219 35224 1619 35240
rect 219 35178 1619 35194
rect 219 35144 231 35178
rect 1607 35144 1619 35178
rect 219 35128 1619 35144
rect 219 35082 1619 35098
rect 219 35048 231 35082
rect 1607 35048 1619 35082
rect 219 35032 1619 35048
rect 219 34986 1619 35002
rect 219 34952 231 34986
rect 1607 34952 1619 34986
rect 219 34936 1619 34952
rect 219 34890 1619 34906
rect 219 34856 231 34890
rect 1607 34856 1619 34890
rect 219 34840 1619 34856
rect 219 34794 1619 34810
rect 219 34760 231 34794
rect 1607 34760 1619 34794
rect 219 34744 1619 34760
rect 219 34698 1619 34714
rect 219 34664 231 34698
rect 1607 34664 1619 34698
rect 219 34648 1619 34664
rect 219 34602 1619 34618
rect 219 34568 231 34602
rect 1607 34568 1619 34602
rect 219 34552 1619 34568
rect 219 34506 1619 34522
rect 219 34472 231 34506
rect 1607 34472 1619 34506
rect 219 34456 1619 34472
rect 219 34410 1619 34426
rect 219 34376 231 34410
rect 1607 34376 1619 34410
rect 219 34360 1619 34376
rect 219 34314 1619 34330
rect 219 34280 231 34314
rect 1607 34280 1619 34314
rect 219 34264 1619 34280
rect 219 34218 1619 34234
rect 219 34184 231 34218
rect 1607 34184 1619 34218
rect 219 34168 1619 34184
rect 219 34122 1619 34138
rect 219 34088 231 34122
rect 1607 34088 1619 34122
rect 219 34072 1619 34088
rect 219 34026 1619 34042
rect 219 33992 231 34026
rect 1607 33992 1619 34026
rect 219 33976 1619 33992
rect 219 33930 1619 33946
rect 219 33896 231 33930
rect 1607 33896 1619 33930
rect 219 33880 1619 33896
rect 219 33834 1619 33850
rect 219 33800 231 33834
rect 1607 33800 1619 33834
rect 219 33784 1619 33800
rect 219 33738 1619 33754
rect 219 33704 231 33738
rect 1607 33704 1619 33738
rect 219 33688 1619 33704
rect 219 33642 1619 33658
rect 219 33608 231 33642
rect 1607 33608 1619 33642
rect 219 33592 1619 33608
rect 219 33546 1619 33562
rect 219 33512 231 33546
rect 1607 33512 1619 33546
rect 219 33496 1619 33512
rect 219 33450 1619 33466
rect 219 33416 231 33450
rect 1607 33416 1619 33450
rect 219 33400 1619 33416
rect 219 33354 1619 33370
rect 219 33320 231 33354
rect 1607 33320 1619 33354
rect 219 33304 1619 33320
rect 219 33258 1619 33274
rect 219 33224 231 33258
rect 1607 33224 1619 33258
rect 219 33208 1619 33224
rect 219 33162 1619 33178
rect 219 33128 231 33162
rect 1607 33128 1619 33162
rect 219 33112 1619 33128
rect 219 33066 1619 33082
rect 219 33032 231 33066
rect 1607 33032 1619 33066
rect 219 33016 1619 33032
rect 219 32970 1619 32986
rect 219 32936 231 32970
rect 1607 32936 1619 32970
rect 219 32920 1619 32936
rect 219 32874 1619 32890
rect 219 32840 231 32874
rect 1607 32840 1619 32874
rect 219 32824 1619 32840
rect 219 32778 1619 32794
rect 219 32744 231 32778
rect 1607 32744 1619 32778
rect 219 32728 1619 32744
rect 219 32682 1619 32698
rect 219 32648 231 32682
rect 1607 32648 1619 32682
rect 219 32632 1619 32648
rect 219 32586 1619 32602
rect 219 32552 231 32586
rect 1607 32552 1619 32586
rect 219 32536 1619 32552
rect 219 32490 1619 32506
rect 219 32456 231 32490
rect 1607 32456 1619 32490
rect 219 32440 1619 32456
rect 219 32394 1619 32410
rect 219 32360 231 32394
rect 1607 32360 1619 32394
rect 219 32344 1619 32360
rect 219 32298 1619 32314
rect 219 32264 231 32298
rect 1607 32264 1619 32298
rect 219 32248 1619 32264
rect 219 32202 1619 32218
rect 219 32168 231 32202
rect 1607 32168 1619 32202
rect 219 32152 1619 32168
rect 219 32106 1619 32122
rect 219 32072 231 32106
rect 1607 32072 1619 32106
rect 219 32056 1619 32072
rect 219 32010 1619 32026
rect 219 31976 231 32010
rect 1607 31976 1619 32010
rect 219 31960 1619 31976
rect 219 31914 1619 31930
rect 219 31880 231 31914
rect 1607 31880 1619 31914
rect 219 31864 1619 31880
rect 219 31818 1619 31834
rect 219 31784 231 31818
rect 1607 31784 1619 31818
rect 219 31768 1619 31784
rect 219 31722 1619 31738
rect 219 31688 231 31722
rect 1607 31688 1619 31722
rect 219 31672 1619 31688
rect 219 31626 1619 31642
rect 219 31592 231 31626
rect 1607 31592 1619 31626
rect 219 31576 1619 31592
rect 219 31530 1619 31546
rect 219 31496 231 31530
rect 1607 31496 1619 31530
rect 219 31480 1619 31496
rect 219 31434 1619 31450
rect 219 31400 231 31434
rect 1607 31400 1619 31434
rect 219 31384 1619 31400
rect 219 31338 1619 31354
rect 219 31304 231 31338
rect 1607 31304 1619 31338
rect 219 31288 1619 31304
rect 219 31242 1619 31258
rect 219 31208 231 31242
rect 1607 31208 1619 31242
rect 219 31192 1619 31208
rect 219 31146 1619 31162
rect 219 31112 231 31146
rect 1607 31112 1619 31146
rect 219 31096 1619 31112
rect 219 31050 1619 31066
rect 219 31016 231 31050
rect 1607 31016 1619 31050
rect 219 31000 1619 31016
rect 219 30954 1619 30970
rect 219 30920 231 30954
rect 1607 30920 1619 30954
rect 219 30904 1619 30920
rect 219 30858 1619 30874
rect 219 30824 231 30858
rect 1607 30824 1619 30858
rect 219 30808 1619 30824
rect 219 30762 1619 30778
rect 219 30728 231 30762
rect 1607 30728 1619 30762
rect 219 30712 1619 30728
rect 219 30666 1619 30682
rect 219 30632 231 30666
rect 1607 30632 1619 30666
rect 219 30616 1619 30632
rect 219 30570 1619 30586
rect 219 30536 231 30570
rect 1607 30536 1619 30570
rect 219 30520 1619 30536
rect 219 30474 1619 30490
rect 219 30440 231 30474
rect 1607 30440 1619 30474
rect 219 30424 1619 30440
rect 219 30378 1619 30394
rect 219 30344 231 30378
rect 1607 30344 1619 30378
rect 219 30328 1619 30344
rect 219 30282 1619 30298
rect 219 30248 231 30282
rect 1607 30248 1619 30282
rect 219 30232 1619 30248
rect 219 30186 1619 30202
rect 219 30152 231 30186
rect 1607 30152 1619 30186
rect 219 30136 1619 30152
rect 219 30090 1619 30106
rect 219 30056 231 30090
rect 1607 30056 1619 30090
rect 219 30040 1619 30056
rect 219 29994 1619 30010
rect 219 29960 231 29994
rect 1607 29960 1619 29994
rect 219 29944 1619 29960
rect 219 29898 1619 29914
rect 219 29864 231 29898
rect 1607 29864 1619 29898
rect 219 29848 1619 29864
rect 219 29802 1619 29818
rect 219 29768 231 29802
rect 1607 29768 1619 29802
rect 219 29752 1619 29768
rect 219 29706 1619 29722
rect 219 29672 231 29706
rect 1607 29672 1619 29706
rect 219 29656 1619 29672
rect 219 29610 1619 29626
rect 219 29576 231 29610
rect 1607 29576 1619 29610
rect 219 29560 1619 29576
rect 219 29514 1619 29530
rect 219 29480 231 29514
rect 1607 29480 1619 29514
rect 219 29464 1619 29480
rect 219 29418 1619 29434
rect 219 29384 231 29418
rect 1607 29384 1619 29418
rect 219 29368 1619 29384
rect 219 29322 1619 29338
rect 219 29288 231 29322
rect 1607 29288 1619 29322
rect 219 29272 1619 29288
rect 219 29226 1619 29242
rect 219 29192 231 29226
rect 1607 29192 1619 29226
rect 219 29176 1619 29192
rect 219 29130 1619 29146
rect 219 29096 231 29130
rect 1607 29096 1619 29130
rect 219 29080 1619 29096
rect 219 29034 1619 29050
rect 219 29000 231 29034
rect 1607 29000 1619 29034
rect 219 28984 1619 29000
rect 219 28938 1619 28954
rect 219 28904 231 28938
rect 1607 28904 1619 28938
rect 219 28888 1619 28904
rect 219 28842 1619 28858
rect 219 28808 231 28842
rect 1607 28808 1619 28842
rect 219 28792 1619 28808
rect 219 28746 1619 28762
rect 219 28712 231 28746
rect 1607 28712 1619 28746
rect 219 28696 1619 28712
rect 219 28650 1619 28666
rect 219 28616 231 28650
rect 1607 28616 1619 28650
rect 219 28600 1619 28616
rect 219 28554 1619 28570
rect 219 28520 231 28554
rect 1607 28520 1619 28554
rect 219 28504 1619 28520
rect 219 28458 1619 28474
rect 219 28424 231 28458
rect 1607 28424 1619 28458
rect 219 28408 1619 28424
rect 219 28362 1619 28378
rect 219 28328 231 28362
rect 1607 28328 1619 28362
rect 219 28312 1619 28328
rect 219 28266 1619 28282
rect 219 28232 231 28266
rect 1607 28232 1619 28266
rect 219 28216 1619 28232
rect 219 28170 1619 28186
rect 219 28136 231 28170
rect 1607 28136 1619 28170
rect 219 28120 1619 28136
rect 219 28074 1619 28090
rect 219 28040 231 28074
rect 1607 28040 1619 28074
rect 219 28024 1619 28040
rect 219 27978 1619 27994
rect 219 27944 231 27978
rect 1607 27944 1619 27978
rect 219 27928 1619 27944
rect 219 27882 1619 27898
rect 219 27848 231 27882
rect 1607 27848 1619 27882
rect 219 27832 1619 27848
rect 219 27786 1619 27802
rect 219 27752 231 27786
rect 1607 27752 1619 27786
rect 219 27736 1619 27752
rect 219 27690 1619 27706
rect 219 27656 231 27690
rect 1607 27656 1619 27690
rect 219 27640 1619 27656
rect 219 27594 1619 27610
rect 219 27560 231 27594
rect 1607 27560 1619 27594
rect 219 27544 1619 27560
rect 219 27498 1619 27514
rect 219 27464 231 27498
rect 1607 27464 1619 27498
rect 219 27448 1619 27464
rect 219 27402 1619 27418
rect 219 27368 231 27402
rect 1607 27368 1619 27402
rect 219 27352 1619 27368
rect 219 27306 1619 27322
rect 219 27272 231 27306
rect 1607 27272 1619 27306
rect 219 27256 1619 27272
rect 219 27210 1619 27226
rect 219 27176 231 27210
rect 1607 27176 1619 27210
rect 219 27160 1619 27176
rect 219 27114 1619 27130
rect 219 27080 231 27114
rect 1607 27080 1619 27114
rect 219 27064 1619 27080
rect 219 27018 1619 27034
rect 219 26984 231 27018
rect 1607 26984 1619 27018
rect 219 26968 1619 26984
rect 219 26922 1619 26938
rect 219 26888 231 26922
rect 1607 26888 1619 26922
rect 219 26872 1619 26888
rect 219 26826 1619 26842
rect 219 26792 231 26826
rect 1607 26792 1619 26826
rect 219 26776 1619 26792
rect 219 26730 1619 26746
rect 219 26696 231 26730
rect 1607 26696 1619 26730
rect 219 26680 1619 26696
rect 219 26634 1619 26650
rect 219 26600 231 26634
rect 1607 26600 1619 26634
rect 219 26584 1619 26600
rect 219 26538 1619 26554
rect 219 26504 231 26538
rect 1607 26504 1619 26538
rect 219 26488 1619 26504
rect 219 26442 1619 26458
rect 219 26408 231 26442
rect 1607 26408 1619 26442
rect 219 26392 1619 26408
rect 219 26346 1619 26362
rect 219 26312 231 26346
rect 1607 26312 1619 26346
rect 219 26296 1619 26312
rect 219 26250 1619 26266
rect 219 26216 231 26250
rect 1607 26216 1619 26250
rect 219 26200 1619 26216
rect 219 26154 1619 26170
rect 219 26120 231 26154
rect 1607 26120 1619 26154
rect 219 26104 1619 26120
rect 219 26058 1619 26074
rect 219 26024 231 26058
rect 1607 26024 1619 26058
rect 219 26008 1619 26024
rect 219 25962 1619 25978
rect 219 25928 231 25962
rect 1607 25928 1619 25962
rect 219 25912 1619 25928
rect 219 25866 1619 25882
rect 219 25832 231 25866
rect 1607 25832 1619 25866
rect 219 25816 1619 25832
rect 219 25770 1619 25786
rect 219 25736 231 25770
rect 1607 25736 1619 25770
rect 219 25720 1619 25736
rect 219 25674 1619 25690
rect 219 25640 231 25674
rect 1607 25640 1619 25674
rect 219 25624 1619 25640
rect 219 25578 1619 25594
rect 219 25544 231 25578
rect 1607 25544 1619 25578
rect 219 25528 1619 25544
rect 219 25482 1619 25498
rect 219 25448 231 25482
rect 1607 25448 1619 25482
rect 219 25432 1619 25448
rect 219 25386 1619 25402
rect 219 25352 231 25386
rect 1607 25352 1619 25386
rect 219 25336 1619 25352
rect 219 25290 1619 25306
rect 219 25256 231 25290
rect 1607 25256 1619 25290
rect 219 25240 1619 25256
rect 219 25194 1619 25210
rect 219 25160 231 25194
rect 1607 25160 1619 25194
rect 219 25144 1619 25160
rect 219 25098 1619 25114
rect 219 25064 231 25098
rect 1607 25064 1619 25098
rect 219 25048 1619 25064
rect 219 25002 1619 25018
rect 219 24968 231 25002
rect 1607 24968 1619 25002
rect 219 24952 1619 24968
rect 219 24906 1619 24922
rect 219 24872 231 24906
rect 1607 24872 1619 24906
rect 219 24856 1619 24872
rect 219 24810 1619 24826
rect 219 24776 231 24810
rect 1607 24776 1619 24810
rect 219 24760 1619 24776
rect 219 24714 1619 24730
rect 219 24680 231 24714
rect 1607 24680 1619 24714
rect 219 24664 1619 24680
rect 219 24618 1619 24634
rect 219 24584 231 24618
rect 1607 24584 1619 24618
rect 219 24568 1619 24584
rect 219 24522 1619 24538
rect 219 24488 231 24522
rect 1607 24488 1619 24522
rect 219 24472 1619 24488
rect 219 24426 1619 24442
rect 219 24392 231 24426
rect 1607 24392 1619 24426
rect 219 24376 1619 24392
rect 219 24330 1619 24346
rect 219 24296 231 24330
rect 1607 24296 1619 24330
rect 219 24280 1619 24296
rect 219 24234 1619 24250
rect 219 24200 231 24234
rect 1607 24200 1619 24234
rect 219 24184 1619 24200
rect 219 24138 1619 24154
rect 219 24104 231 24138
rect 1607 24104 1619 24138
rect 219 24088 1619 24104
rect 219 24042 1619 24058
rect 219 24008 231 24042
rect 1607 24008 1619 24042
rect 219 23992 1619 24008
rect 219 23946 1619 23962
rect 219 23912 231 23946
rect 1607 23912 1619 23946
rect 219 23896 1619 23912
rect 219 23850 1619 23866
rect 219 23816 231 23850
rect 1607 23816 1619 23850
rect 219 23800 1619 23816
rect 219 23754 1619 23770
rect 219 23720 231 23754
rect 1607 23720 1619 23754
rect 219 23704 1619 23720
rect 219 23658 1619 23674
rect 219 23624 231 23658
rect 1607 23624 1619 23658
rect 219 23608 1619 23624
rect 219 23562 1619 23578
rect 219 23528 231 23562
rect 1607 23528 1619 23562
rect 219 23512 1619 23528
rect 219 23466 1619 23482
rect 219 23432 231 23466
rect 1607 23432 1619 23466
rect 219 23416 1619 23432
rect 219 23370 1619 23386
rect 219 23336 231 23370
rect 1607 23336 1619 23370
rect 219 23320 1619 23336
rect 219 23274 1619 23290
rect 219 23240 231 23274
rect 1607 23240 1619 23274
rect 219 23224 1619 23240
rect 219 23178 1619 23194
rect 219 23144 231 23178
rect 1607 23144 1619 23178
rect 219 23128 1619 23144
rect 219 23082 1619 23098
rect 219 23048 231 23082
rect 1607 23048 1619 23082
rect 219 23036 1619 23048
rect 219 21704 1619 21716
rect 219 21670 231 21704
rect 1607 21670 1619 21704
rect 219 21654 1619 21670
rect 219 21608 1619 21624
rect 219 21574 231 21608
rect 1607 21574 1619 21608
rect 219 21558 1619 21574
rect 219 21512 1619 21528
rect 219 21478 231 21512
rect 1607 21478 1619 21512
rect 219 21462 1619 21478
rect 219 21416 1619 21432
rect 219 21382 231 21416
rect 1607 21382 1619 21416
rect 219 21366 1619 21382
rect 219 21320 1619 21336
rect 219 21286 231 21320
rect 1607 21286 1619 21320
rect 219 21270 1619 21286
rect 219 21224 1619 21240
rect 219 21190 231 21224
rect 1607 21190 1619 21224
rect 219 21174 1619 21190
rect 219 21128 1619 21144
rect 219 21094 231 21128
rect 1607 21094 1619 21128
rect 219 21078 1619 21094
rect 219 21032 1619 21048
rect 219 20998 231 21032
rect 1607 20998 1619 21032
rect 219 20982 1619 20998
rect 219 20936 1619 20952
rect 219 20902 231 20936
rect 1607 20902 1619 20936
rect 219 20886 1619 20902
rect 219 20840 1619 20856
rect 219 20806 231 20840
rect 1607 20806 1619 20840
rect 219 20790 1619 20806
rect 219 20744 1619 20760
rect 219 20710 231 20744
rect 1607 20710 1619 20744
rect 219 20694 1619 20710
rect 219 20648 1619 20664
rect 219 20614 231 20648
rect 1607 20614 1619 20648
rect 219 20598 1619 20614
rect 219 20552 1619 20568
rect 219 20518 231 20552
rect 1607 20518 1619 20552
rect 219 20502 1619 20518
rect 219 20456 1619 20472
rect 219 20422 231 20456
rect 1607 20422 1619 20456
rect 219 20406 1619 20422
rect 219 20360 1619 20376
rect 219 20326 231 20360
rect 1607 20326 1619 20360
rect 219 20310 1619 20326
rect 219 20264 1619 20280
rect 219 20230 231 20264
rect 1607 20230 1619 20264
rect 219 20214 1619 20230
rect 219 20168 1619 20184
rect 219 20134 231 20168
rect 1607 20134 1619 20168
rect 219 20118 1619 20134
rect 219 20072 1619 20088
rect 219 20038 231 20072
rect 1607 20038 1619 20072
rect 219 20022 1619 20038
rect 219 19976 1619 19992
rect 219 19942 231 19976
rect 1607 19942 1619 19976
rect 219 19926 1619 19942
rect 219 19880 1619 19896
rect 219 19846 231 19880
rect 1607 19846 1619 19880
rect 219 19830 1619 19846
rect 219 19784 1619 19800
rect 219 19750 231 19784
rect 1607 19750 1619 19784
rect 219 19734 1619 19750
rect 219 19688 1619 19704
rect 219 19654 231 19688
rect 1607 19654 1619 19688
rect 219 19638 1619 19654
rect 219 19592 1619 19608
rect 219 19558 231 19592
rect 1607 19558 1619 19592
rect 219 19542 1619 19558
rect 219 19496 1619 19512
rect 219 19462 231 19496
rect 1607 19462 1619 19496
rect 219 19446 1619 19462
rect 219 19400 1619 19416
rect 219 19366 231 19400
rect 1607 19366 1619 19400
rect 219 19350 1619 19366
rect 219 19304 1619 19320
rect 219 19270 231 19304
rect 1607 19270 1619 19304
rect 219 19254 1619 19270
rect 219 19208 1619 19224
rect 219 19174 231 19208
rect 1607 19174 1619 19208
rect 219 19158 1619 19174
rect 219 19112 1619 19128
rect 219 19078 231 19112
rect 1607 19078 1619 19112
rect 219 19062 1619 19078
rect 219 19016 1619 19032
rect 219 18982 231 19016
rect 1607 18982 1619 19016
rect 219 18966 1619 18982
rect 219 18920 1619 18936
rect 219 18886 231 18920
rect 1607 18886 1619 18920
rect 219 18870 1619 18886
rect 219 18824 1619 18840
rect 219 18790 231 18824
rect 1607 18790 1619 18824
rect 219 18774 1619 18790
rect 219 18728 1619 18744
rect 219 18694 231 18728
rect 1607 18694 1619 18728
rect 219 18678 1619 18694
rect 219 18632 1619 18648
rect 219 18598 231 18632
rect 1607 18598 1619 18632
rect 219 18582 1619 18598
rect 219 18536 1619 18552
rect 219 18502 231 18536
rect 1607 18502 1619 18536
rect 219 18486 1619 18502
rect 219 18440 1619 18456
rect 219 18406 231 18440
rect 1607 18406 1619 18440
rect 219 18390 1619 18406
rect 219 18344 1619 18360
rect 219 18310 231 18344
rect 1607 18310 1619 18344
rect 219 18294 1619 18310
rect 219 18248 1619 18264
rect 219 18214 231 18248
rect 1607 18214 1619 18248
rect 219 18198 1619 18214
rect 219 18152 1619 18168
rect 219 18118 231 18152
rect 1607 18118 1619 18152
rect 219 18102 1619 18118
rect 219 18056 1619 18072
rect 219 18022 231 18056
rect 1607 18022 1619 18056
rect 219 18006 1619 18022
rect 219 17960 1619 17976
rect 219 17926 231 17960
rect 1607 17926 1619 17960
rect 219 17910 1619 17926
rect 219 17864 1619 17880
rect 219 17830 231 17864
rect 1607 17830 1619 17864
rect 219 17814 1619 17830
rect 219 17768 1619 17784
rect 219 17734 231 17768
rect 1607 17734 1619 17768
rect 219 17718 1619 17734
rect 219 17672 1619 17688
rect 219 17638 231 17672
rect 1607 17638 1619 17672
rect 219 17622 1619 17638
rect 219 17576 1619 17592
rect 219 17542 231 17576
rect 1607 17542 1619 17576
rect 219 17526 1619 17542
rect 219 17480 1619 17496
rect 219 17446 231 17480
rect 1607 17446 1619 17480
rect 219 17430 1619 17446
rect 219 17384 1619 17400
rect 219 17350 231 17384
rect 1607 17350 1619 17384
rect 219 17334 1619 17350
rect 219 17288 1619 17304
rect 219 17254 231 17288
rect 1607 17254 1619 17288
rect 219 17238 1619 17254
rect 219 17192 1619 17208
rect 219 17158 231 17192
rect 1607 17158 1619 17192
rect 219 17142 1619 17158
rect 219 17096 1619 17112
rect 219 17062 231 17096
rect 1607 17062 1619 17096
rect 219 17046 1619 17062
rect 219 17000 1619 17016
rect 219 16966 231 17000
rect 1607 16966 1619 17000
rect 219 16950 1619 16966
rect 219 16904 1619 16920
rect 219 16870 231 16904
rect 1607 16870 1619 16904
rect 219 16854 1619 16870
rect 219 16808 1619 16824
rect 219 16774 231 16808
rect 1607 16774 1619 16808
rect 219 16758 1619 16774
rect 219 16712 1619 16728
rect 219 16678 231 16712
rect 1607 16678 1619 16712
rect 219 16662 1619 16678
rect 219 16616 1619 16632
rect 219 16582 231 16616
rect 1607 16582 1619 16616
rect 219 16566 1619 16582
rect 219 16520 1619 16536
rect 219 16486 231 16520
rect 1607 16486 1619 16520
rect 219 16470 1619 16486
rect 219 16424 1619 16440
rect 219 16390 231 16424
rect 1607 16390 1619 16424
rect 219 16374 1619 16390
rect 219 16328 1619 16344
rect 219 16294 231 16328
rect 1607 16294 1619 16328
rect 219 16278 1619 16294
rect 219 16232 1619 16248
rect 219 16198 231 16232
rect 1607 16198 1619 16232
rect 219 16182 1619 16198
rect 219 16136 1619 16152
rect 219 16102 231 16136
rect 1607 16102 1619 16136
rect 219 16086 1619 16102
rect 219 16040 1619 16056
rect 219 16006 231 16040
rect 1607 16006 1619 16040
rect 219 15990 1619 16006
rect 219 15944 1619 15960
rect 219 15910 231 15944
rect 1607 15910 1619 15944
rect 219 15894 1619 15910
rect 219 15848 1619 15864
rect 219 15814 231 15848
rect 1607 15814 1619 15848
rect 219 15798 1619 15814
rect 219 15752 1619 15768
rect 219 15718 231 15752
rect 1607 15718 1619 15752
rect 219 15702 1619 15718
rect 219 15656 1619 15672
rect 219 15622 231 15656
rect 1607 15622 1619 15656
rect 219 15606 1619 15622
rect 219 15560 1619 15576
rect 219 15526 231 15560
rect 1607 15526 1619 15560
rect 219 15510 1619 15526
rect 219 15464 1619 15480
rect 219 15430 231 15464
rect 1607 15430 1619 15464
rect 219 15414 1619 15430
rect 219 15368 1619 15384
rect 219 15334 231 15368
rect 1607 15334 1619 15368
rect 219 15318 1619 15334
rect 219 15272 1619 15288
rect 219 15238 231 15272
rect 1607 15238 1619 15272
rect 219 15222 1619 15238
rect 219 15176 1619 15192
rect 219 15142 231 15176
rect 1607 15142 1619 15176
rect 219 15126 1619 15142
rect 219 15080 1619 15096
rect 219 15046 231 15080
rect 1607 15046 1619 15080
rect 219 15030 1619 15046
rect 219 14984 1619 15000
rect 219 14950 231 14984
rect 1607 14950 1619 14984
rect 219 14934 1619 14950
rect 219 14888 1619 14904
rect 219 14854 231 14888
rect 1607 14854 1619 14888
rect 219 14838 1619 14854
rect 219 14792 1619 14808
rect 219 14758 231 14792
rect 1607 14758 1619 14792
rect 219 14742 1619 14758
rect 219 14696 1619 14712
rect 219 14662 231 14696
rect 1607 14662 1619 14696
rect 219 14646 1619 14662
rect 219 14600 1619 14616
rect 219 14566 231 14600
rect 1607 14566 1619 14600
rect 219 14550 1619 14566
rect 219 14504 1619 14520
rect 219 14470 231 14504
rect 1607 14470 1619 14504
rect 219 14454 1619 14470
rect 219 14408 1619 14424
rect 219 14374 231 14408
rect 1607 14374 1619 14408
rect 219 14358 1619 14374
rect 219 14312 1619 14328
rect 219 14278 231 14312
rect 1607 14278 1619 14312
rect 219 14262 1619 14278
rect 219 14216 1619 14232
rect 219 14182 231 14216
rect 1607 14182 1619 14216
rect 219 14166 1619 14182
rect 219 14120 1619 14136
rect 219 14086 231 14120
rect 1607 14086 1619 14120
rect 219 14070 1619 14086
rect 219 14024 1619 14040
rect 219 13990 231 14024
rect 1607 13990 1619 14024
rect 219 13974 1619 13990
rect 219 13928 1619 13944
rect 219 13894 231 13928
rect 1607 13894 1619 13928
rect 219 13878 1619 13894
rect 219 13832 1619 13848
rect 219 13798 231 13832
rect 1607 13798 1619 13832
rect 219 13782 1619 13798
rect 219 13736 1619 13752
rect 219 13702 231 13736
rect 1607 13702 1619 13736
rect 219 13686 1619 13702
rect 219 13640 1619 13656
rect 219 13606 231 13640
rect 1607 13606 1619 13640
rect 219 13590 1619 13606
rect 219 13544 1619 13560
rect 219 13510 231 13544
rect 1607 13510 1619 13544
rect 219 13494 1619 13510
rect 219 13448 1619 13464
rect 219 13414 231 13448
rect 1607 13414 1619 13448
rect 219 13398 1619 13414
rect 219 13352 1619 13368
rect 219 13318 231 13352
rect 1607 13318 1619 13352
rect 219 13302 1619 13318
rect 219 13256 1619 13272
rect 219 13222 231 13256
rect 1607 13222 1619 13256
rect 219 13206 1619 13222
rect 219 13160 1619 13176
rect 219 13126 231 13160
rect 1607 13126 1619 13160
rect 219 13110 1619 13126
rect 219 13064 1619 13080
rect 219 13030 231 13064
rect 1607 13030 1619 13064
rect 219 13014 1619 13030
rect 219 12968 1619 12984
rect 219 12934 231 12968
rect 1607 12934 1619 12968
rect 219 12918 1619 12934
rect 219 12872 1619 12888
rect 219 12838 231 12872
rect 1607 12838 1619 12872
rect 219 12822 1619 12838
rect 219 12776 1619 12792
rect 219 12742 231 12776
rect 1607 12742 1619 12776
rect 219 12726 1619 12742
rect 219 12680 1619 12696
rect 219 12646 231 12680
rect 1607 12646 1619 12680
rect 219 12630 1619 12646
rect 219 12584 1619 12600
rect 219 12550 231 12584
rect 1607 12550 1619 12584
rect 219 12534 1619 12550
rect 219 12488 1619 12504
rect 219 12454 231 12488
rect 1607 12454 1619 12488
rect 219 12438 1619 12454
rect 219 12392 1619 12408
rect 219 12358 231 12392
rect 1607 12358 1619 12392
rect 219 12342 1619 12358
rect 219 12296 1619 12312
rect 219 12262 231 12296
rect 1607 12262 1619 12296
rect 219 12246 1619 12262
rect 219 12200 1619 12216
rect 219 12166 231 12200
rect 1607 12166 1619 12200
rect 219 12150 1619 12166
rect 219 12104 1619 12120
rect 219 12070 231 12104
rect 1607 12070 1619 12104
rect 219 12054 1619 12070
rect 219 12008 1619 12024
rect 219 11974 231 12008
rect 1607 11974 1619 12008
rect 219 11958 1619 11974
rect 219 11912 1619 11928
rect 219 11878 231 11912
rect 1607 11878 1619 11912
rect 219 11862 1619 11878
rect 219 11816 1619 11832
rect 219 11782 231 11816
rect 1607 11782 1619 11816
rect 219 11766 1619 11782
rect 219 11720 1619 11736
rect 219 11686 231 11720
rect 1607 11686 1619 11720
rect 219 11670 1619 11686
rect 219 11624 1619 11640
rect 219 11590 231 11624
rect 1607 11590 1619 11624
rect 219 11574 1619 11590
rect 219 11528 1619 11544
rect 219 11494 231 11528
rect 1607 11494 1619 11528
rect 219 11478 1619 11494
rect 219 11432 1619 11448
rect 219 11398 231 11432
rect 1607 11398 1619 11432
rect 219 11382 1619 11398
rect 219 11336 1619 11352
rect 219 11302 231 11336
rect 1607 11302 1619 11336
rect 219 11286 1619 11302
rect 219 11240 1619 11256
rect 219 11206 231 11240
rect 1607 11206 1619 11240
rect 219 11190 1619 11206
rect 219 11144 1619 11160
rect 219 11110 231 11144
rect 1607 11110 1619 11144
rect 219 11094 1619 11110
rect 219 11048 1619 11064
rect 219 11014 231 11048
rect 1607 11014 1619 11048
rect 219 10998 1619 11014
rect 219 10952 1619 10968
rect 219 10918 231 10952
rect 1607 10918 1619 10952
rect 219 10902 1619 10918
rect 219 10856 1619 10872
rect 219 10822 231 10856
rect 1607 10822 1619 10856
rect 219 10806 1619 10822
rect 219 10760 1619 10776
rect 219 10726 231 10760
rect 1607 10726 1619 10760
rect 219 10710 1619 10726
rect 219 10664 1619 10680
rect 219 10630 231 10664
rect 1607 10630 1619 10664
rect 219 10614 1619 10630
rect 219 10568 1619 10584
rect 219 10534 231 10568
rect 1607 10534 1619 10568
rect 219 10518 1619 10534
rect 219 10472 1619 10488
rect 219 10438 231 10472
rect 1607 10438 1619 10472
rect 219 10422 1619 10438
rect 219 10376 1619 10392
rect 219 10342 231 10376
rect 1607 10342 1619 10376
rect 219 10326 1619 10342
rect 219 10280 1619 10296
rect 219 10246 231 10280
rect 1607 10246 1619 10280
rect 219 10230 1619 10246
rect 219 10184 1619 10200
rect 219 10150 231 10184
rect 1607 10150 1619 10184
rect 219 10134 1619 10150
rect 219 10088 1619 10104
rect 219 10054 231 10088
rect 1607 10054 1619 10088
rect 219 10038 1619 10054
rect 219 9992 1619 10008
rect 219 9958 231 9992
rect 1607 9958 1619 9992
rect 219 9942 1619 9958
rect 219 9896 1619 9912
rect 219 9862 231 9896
rect 1607 9862 1619 9896
rect 219 9846 1619 9862
rect 219 9800 1619 9816
rect 219 9766 231 9800
rect 1607 9766 1619 9800
rect 219 9750 1619 9766
rect 219 9704 1619 9720
rect 219 9670 231 9704
rect 1607 9670 1619 9704
rect 219 9654 1619 9670
rect 219 9608 1619 9624
rect 219 9574 231 9608
rect 1607 9574 1619 9608
rect 219 9558 1619 9574
rect 219 9512 1619 9528
rect 219 9478 231 9512
rect 1607 9478 1619 9512
rect 219 9462 1619 9478
rect 219 9416 1619 9432
rect 219 9382 231 9416
rect 1607 9382 1619 9416
rect 219 9366 1619 9382
rect 219 9320 1619 9336
rect 219 9286 231 9320
rect 1607 9286 1619 9320
rect 219 9270 1619 9286
rect 219 9224 1619 9240
rect 219 9190 231 9224
rect 1607 9190 1619 9224
rect 219 9174 1619 9190
rect 219 9128 1619 9144
rect 219 9094 231 9128
rect 1607 9094 1619 9128
rect 219 9078 1619 9094
rect 219 9032 1619 9048
rect 219 8998 231 9032
rect 1607 8998 1619 9032
rect 219 8982 1619 8998
rect 219 8936 1619 8952
rect 219 8902 231 8936
rect 1607 8902 1619 8936
rect 219 8886 1619 8902
rect 219 8840 1619 8856
rect 219 8806 231 8840
rect 1607 8806 1619 8840
rect 219 8790 1619 8806
rect 219 8744 1619 8760
rect 219 8710 231 8744
rect 1607 8710 1619 8744
rect 219 8694 1619 8710
rect 219 8648 1619 8664
rect 219 8614 231 8648
rect 1607 8614 1619 8648
rect 219 8598 1619 8614
rect 219 8552 1619 8568
rect 219 8518 231 8552
rect 1607 8518 1619 8552
rect 219 8502 1619 8518
rect 219 8456 1619 8472
rect 219 8422 231 8456
rect 1607 8422 1619 8456
rect 219 8406 1619 8422
rect 219 8360 1619 8376
rect 219 8326 231 8360
rect 1607 8326 1619 8360
rect 219 8310 1619 8326
rect 219 8264 1619 8280
rect 219 8230 231 8264
rect 1607 8230 1619 8264
rect 219 8214 1619 8230
rect 219 8168 1619 8184
rect 219 8134 231 8168
rect 1607 8134 1619 8168
rect 219 8118 1619 8134
rect 219 8072 1619 8088
rect 219 8038 231 8072
rect 1607 8038 1619 8072
rect 219 8022 1619 8038
rect 219 7976 1619 7992
rect 219 7942 231 7976
rect 1607 7942 1619 7976
rect 219 7926 1619 7942
rect 219 7880 1619 7896
rect 219 7846 231 7880
rect 1607 7846 1619 7880
rect 219 7830 1619 7846
rect 219 7784 1619 7800
rect 219 7750 231 7784
rect 1607 7750 1619 7784
rect 219 7734 1619 7750
rect 219 7688 1619 7704
rect 219 7654 231 7688
rect 1607 7654 1619 7688
rect 219 7638 1619 7654
rect 219 7592 1619 7608
rect 219 7558 231 7592
rect 1607 7558 1619 7592
rect 219 7542 1619 7558
rect 219 7496 1619 7512
rect 219 7462 231 7496
rect 1607 7462 1619 7496
rect 219 7446 1619 7462
rect 219 7400 1619 7416
rect 219 7366 231 7400
rect 1607 7366 1619 7400
rect 219 7350 1619 7366
rect 219 7304 1619 7320
rect 219 7270 231 7304
rect 1607 7270 1619 7304
rect 219 7254 1619 7270
rect 219 7208 1619 7224
rect 219 7174 231 7208
rect 1607 7174 1619 7208
rect 219 7158 1619 7174
rect 219 7112 1619 7128
rect 219 7078 231 7112
rect 1607 7078 1619 7112
rect 219 7062 1619 7078
rect 219 7016 1619 7032
rect 219 6982 231 7016
rect 1607 6982 1619 7016
rect 219 6966 1619 6982
rect 219 6920 1619 6936
rect 219 6886 231 6920
rect 1607 6886 1619 6920
rect 219 6870 1619 6886
rect 219 6824 1619 6840
rect 219 6790 231 6824
rect 1607 6790 1619 6824
rect 219 6774 1619 6790
rect 219 6728 1619 6744
rect 219 6694 231 6728
rect 1607 6694 1619 6728
rect 219 6678 1619 6694
rect 219 6632 1619 6648
rect 219 6598 231 6632
rect 1607 6598 1619 6632
rect 219 6582 1619 6598
rect 219 6536 1619 6552
rect 219 6502 231 6536
rect 1607 6502 1619 6536
rect 219 6486 1619 6502
rect 219 6440 1619 6456
rect 219 6406 231 6440
rect 1607 6406 1619 6440
rect 219 6390 1619 6406
rect 219 6344 1619 6360
rect 219 6310 231 6344
rect 1607 6310 1619 6344
rect 219 6294 1619 6310
rect 219 6248 1619 6264
rect 219 6214 231 6248
rect 1607 6214 1619 6248
rect 219 6198 1619 6214
rect 219 6152 1619 6168
rect 219 6118 231 6152
rect 1607 6118 1619 6152
rect 219 6102 1619 6118
rect 219 6056 1619 6072
rect 219 6022 231 6056
rect 1607 6022 1619 6056
rect 219 6006 1619 6022
rect 219 5960 1619 5976
rect 219 5926 231 5960
rect 1607 5926 1619 5960
rect 219 5910 1619 5926
rect 219 5864 1619 5880
rect 219 5830 231 5864
rect 1607 5830 1619 5864
rect 219 5814 1619 5830
rect 219 5768 1619 5784
rect 219 5734 231 5768
rect 1607 5734 1619 5768
rect 219 5718 1619 5734
rect 219 5672 1619 5688
rect 219 5638 231 5672
rect 1607 5638 1619 5672
rect 219 5622 1619 5638
rect 219 5576 1619 5592
rect 219 5542 231 5576
rect 1607 5542 1619 5576
rect 219 5526 1619 5542
rect 219 5480 1619 5496
rect 219 5446 231 5480
rect 1607 5446 1619 5480
rect 219 5430 1619 5446
rect 219 5384 1619 5400
rect 219 5350 231 5384
rect 1607 5350 1619 5384
rect 219 5334 1619 5350
rect 219 5288 1619 5304
rect 219 5254 231 5288
rect 1607 5254 1619 5288
rect 219 5238 1619 5254
rect 219 5192 1619 5208
rect 219 5158 231 5192
rect 1607 5158 1619 5192
rect 219 5142 1619 5158
rect 219 5096 1619 5112
rect 219 5062 231 5096
rect 1607 5062 1619 5096
rect 219 5046 1619 5062
rect 219 5000 1619 5016
rect 219 4966 231 5000
rect 1607 4966 1619 5000
rect 219 4950 1619 4966
rect 219 4904 1619 4920
rect 219 4870 231 4904
rect 1607 4870 1619 4904
rect 219 4854 1619 4870
rect 219 4808 1619 4824
rect 219 4774 231 4808
rect 1607 4774 1619 4808
rect 219 4758 1619 4774
rect 219 4712 1619 4728
rect 219 4678 231 4712
rect 1607 4678 1619 4712
rect 219 4662 1619 4678
rect 219 4616 1619 4632
rect 219 4582 231 4616
rect 1607 4582 1619 4616
rect 219 4566 1619 4582
rect 219 4520 1619 4536
rect 219 4486 231 4520
rect 1607 4486 1619 4520
rect 219 4470 1619 4486
rect 219 4424 1619 4440
rect 219 4390 231 4424
rect 1607 4390 1619 4424
rect 219 4374 1619 4390
rect 219 4328 1619 4344
rect 219 4294 231 4328
rect 1607 4294 1619 4328
rect 219 4278 1619 4294
rect 219 4232 1619 4248
rect 219 4198 231 4232
rect 1607 4198 1619 4232
rect 219 4182 1619 4198
rect 219 4136 1619 4152
rect 219 4102 231 4136
rect 1607 4102 1619 4136
rect 219 4086 1619 4102
rect 219 4040 1619 4056
rect 219 4006 231 4040
rect 1607 4006 1619 4040
rect 219 3990 1619 4006
rect 219 3944 1619 3960
rect 219 3910 231 3944
rect 1607 3910 1619 3944
rect 219 3894 1619 3910
rect 219 3848 1619 3864
rect 219 3814 231 3848
rect 1607 3814 1619 3848
rect 219 3798 1619 3814
rect 219 3752 1619 3768
rect 219 3718 231 3752
rect 1607 3718 1619 3752
rect 219 3702 1619 3718
rect 219 3656 1619 3672
rect 219 3622 231 3656
rect 1607 3622 1619 3656
rect 219 3606 1619 3622
rect 219 3560 1619 3576
rect 219 3526 231 3560
rect 1607 3526 1619 3560
rect 219 3510 1619 3526
rect 219 3464 1619 3480
rect 219 3430 231 3464
rect 1607 3430 1619 3464
rect 219 3414 1619 3430
rect 219 3368 1619 3384
rect 219 3334 231 3368
rect 1607 3334 1619 3368
rect 219 3318 1619 3334
rect 219 3272 1619 3288
rect 219 3238 231 3272
rect 1607 3238 1619 3272
rect 219 3222 1619 3238
rect 219 3176 1619 3192
rect 219 3142 231 3176
rect 1607 3142 1619 3176
rect 219 3126 1619 3142
rect 219 3080 1619 3096
rect 219 3046 231 3080
rect 1607 3046 1619 3080
rect 219 3030 1619 3046
rect 219 2984 1619 3000
rect 219 2950 231 2984
rect 1607 2950 1619 2984
rect 219 2934 1619 2950
rect 219 2888 1619 2904
rect 219 2854 231 2888
rect 1607 2854 1619 2888
rect 219 2838 1619 2854
rect 219 2792 1619 2808
rect 219 2758 231 2792
rect 1607 2758 1619 2792
rect 219 2742 1619 2758
rect 219 2696 1619 2712
rect 219 2662 231 2696
rect 1607 2662 1619 2696
rect 219 2646 1619 2662
rect 219 2600 1619 2616
rect 219 2566 231 2600
rect 1607 2566 1619 2600
rect 219 2550 1619 2566
rect 219 2504 1619 2520
rect 219 2470 231 2504
rect 1607 2470 1619 2504
rect 219 2454 1619 2470
rect 219 2408 1619 2424
rect 219 2374 231 2408
rect 1607 2374 1619 2408
rect 219 2358 1619 2374
rect 219 2312 1619 2328
rect 219 2278 231 2312
rect 1607 2278 1619 2312
rect 219 2262 1619 2278
rect 219 2216 1619 2232
rect 219 2182 231 2216
rect 1607 2182 1619 2216
rect 219 2166 1619 2182
rect 219 2120 1619 2136
rect 219 2086 231 2120
rect 1607 2086 1619 2120
rect 219 2070 1619 2086
rect 219 2024 1619 2040
rect 219 1990 231 2024
rect 1607 1990 1619 2024
rect 219 1974 1619 1990
rect 219 1928 1619 1944
rect 219 1894 231 1928
rect 1607 1894 1619 1928
rect 219 1878 1619 1894
rect 219 1832 1619 1848
rect 219 1798 231 1832
rect 1607 1798 1619 1832
rect 219 1782 1619 1798
rect 219 1736 1619 1752
rect 219 1702 231 1736
rect 1607 1702 1619 1736
rect 219 1686 1619 1702
rect 219 1640 1619 1656
rect 219 1606 231 1640
rect 1607 1606 1619 1640
rect 219 1590 1619 1606
rect 219 1544 1619 1560
rect 219 1510 231 1544
rect 1607 1510 1619 1544
rect 219 1494 1619 1510
rect 219 1448 1619 1464
rect 219 1414 231 1448
rect 1607 1414 1619 1448
rect 219 1398 1619 1414
rect 219 1352 1619 1368
rect 219 1318 231 1352
rect 1607 1318 1619 1352
rect 219 1302 1619 1318
rect 219 1256 1619 1272
rect 219 1222 231 1256
rect 1607 1222 1619 1256
rect 219 1206 1619 1222
rect 219 1160 1619 1176
rect 219 1126 231 1160
rect 1607 1126 1619 1160
rect 219 1110 1619 1126
rect 219 1064 1619 1080
rect 219 1030 231 1064
rect 1607 1030 1619 1064
rect 219 1014 1619 1030
rect 219 968 1619 984
rect 219 934 231 968
rect 1607 934 1619 968
rect 219 918 1619 934
rect 219 872 1619 888
rect 219 838 231 872
rect 1607 838 1619 872
rect 219 822 1619 838
rect 219 776 1619 792
rect 219 742 231 776
rect 1607 742 1619 776
rect 219 726 1619 742
rect 219 680 1619 696
rect 219 646 231 680
rect 1607 646 1619 680
rect 219 630 1619 646
rect 219 584 1619 600
rect 219 550 231 584
rect 1607 550 1619 584
rect 219 538 1619 550
<< pdiffc >>
rect 231 44168 1607 44202
rect 231 44072 1607 44106
rect 231 43976 1607 44010
rect 231 43880 1607 43914
rect 231 43784 1607 43818
rect 231 43688 1607 43722
rect 231 43592 1607 43626
rect 231 43496 1607 43530
rect 231 43400 1607 43434
rect 231 43304 1607 43338
rect 231 43208 1607 43242
rect 231 43112 1607 43146
rect 231 43016 1607 43050
rect 231 42920 1607 42954
rect 231 42824 1607 42858
rect 231 42728 1607 42762
rect 231 42632 1607 42666
rect 231 42536 1607 42570
rect 231 42440 1607 42474
rect 231 42344 1607 42378
rect 231 42248 1607 42282
rect 231 42152 1607 42186
rect 231 42056 1607 42090
rect 231 41960 1607 41994
rect 231 41864 1607 41898
rect 231 41768 1607 41802
rect 231 41672 1607 41706
rect 231 41576 1607 41610
rect 231 41480 1607 41514
rect 231 41384 1607 41418
rect 231 41288 1607 41322
rect 231 41192 1607 41226
rect 231 41096 1607 41130
rect 231 41000 1607 41034
rect 231 40904 1607 40938
rect 231 40808 1607 40842
rect 231 40712 1607 40746
rect 231 40616 1607 40650
rect 231 40520 1607 40554
rect 231 40424 1607 40458
rect 231 40328 1607 40362
rect 231 40232 1607 40266
rect 231 40136 1607 40170
rect 231 40040 1607 40074
rect 231 39944 1607 39978
rect 231 39848 1607 39882
rect 231 39752 1607 39786
rect 231 39656 1607 39690
rect 231 39560 1607 39594
rect 231 39464 1607 39498
rect 231 39368 1607 39402
rect 231 39272 1607 39306
rect 231 39176 1607 39210
rect 231 39080 1607 39114
rect 231 38984 1607 39018
rect 231 38888 1607 38922
rect 231 38792 1607 38826
rect 231 38696 1607 38730
rect 231 38600 1607 38634
rect 231 38504 1607 38538
rect 231 38408 1607 38442
rect 231 38312 1607 38346
rect 231 38216 1607 38250
rect 231 38120 1607 38154
rect 231 38024 1607 38058
rect 231 37928 1607 37962
rect 231 37832 1607 37866
rect 231 37736 1607 37770
rect 231 37640 1607 37674
rect 231 37544 1607 37578
rect 231 37448 1607 37482
rect 231 37352 1607 37386
rect 231 37256 1607 37290
rect 231 37160 1607 37194
rect 231 37064 1607 37098
rect 231 36968 1607 37002
rect 231 36872 1607 36906
rect 231 36776 1607 36810
rect 231 36680 1607 36714
rect 231 36584 1607 36618
rect 231 36488 1607 36522
rect 231 36392 1607 36426
rect 231 36296 1607 36330
rect 231 36200 1607 36234
rect 231 36104 1607 36138
rect 231 36008 1607 36042
rect 231 35912 1607 35946
rect 231 35816 1607 35850
rect 231 35720 1607 35754
rect 231 35624 1607 35658
rect 231 35528 1607 35562
rect 231 35432 1607 35466
rect 231 35336 1607 35370
rect 231 35240 1607 35274
rect 231 35144 1607 35178
rect 231 35048 1607 35082
rect 231 34952 1607 34986
rect 231 34856 1607 34890
rect 231 34760 1607 34794
rect 231 34664 1607 34698
rect 231 34568 1607 34602
rect 231 34472 1607 34506
rect 231 34376 1607 34410
rect 231 34280 1607 34314
rect 231 34184 1607 34218
rect 231 34088 1607 34122
rect 231 33992 1607 34026
rect 231 33896 1607 33930
rect 231 33800 1607 33834
rect 231 33704 1607 33738
rect 231 33608 1607 33642
rect 231 33512 1607 33546
rect 231 33416 1607 33450
rect 231 33320 1607 33354
rect 231 33224 1607 33258
rect 231 33128 1607 33162
rect 231 33032 1607 33066
rect 231 32936 1607 32970
rect 231 32840 1607 32874
rect 231 32744 1607 32778
rect 231 32648 1607 32682
rect 231 32552 1607 32586
rect 231 32456 1607 32490
rect 231 32360 1607 32394
rect 231 32264 1607 32298
rect 231 32168 1607 32202
rect 231 32072 1607 32106
rect 231 31976 1607 32010
rect 231 31880 1607 31914
rect 231 31784 1607 31818
rect 231 31688 1607 31722
rect 231 31592 1607 31626
rect 231 31496 1607 31530
rect 231 31400 1607 31434
rect 231 31304 1607 31338
rect 231 31208 1607 31242
rect 231 31112 1607 31146
rect 231 31016 1607 31050
rect 231 30920 1607 30954
rect 231 30824 1607 30858
rect 231 30728 1607 30762
rect 231 30632 1607 30666
rect 231 30536 1607 30570
rect 231 30440 1607 30474
rect 231 30344 1607 30378
rect 231 30248 1607 30282
rect 231 30152 1607 30186
rect 231 30056 1607 30090
rect 231 29960 1607 29994
rect 231 29864 1607 29898
rect 231 29768 1607 29802
rect 231 29672 1607 29706
rect 231 29576 1607 29610
rect 231 29480 1607 29514
rect 231 29384 1607 29418
rect 231 29288 1607 29322
rect 231 29192 1607 29226
rect 231 29096 1607 29130
rect 231 29000 1607 29034
rect 231 28904 1607 28938
rect 231 28808 1607 28842
rect 231 28712 1607 28746
rect 231 28616 1607 28650
rect 231 28520 1607 28554
rect 231 28424 1607 28458
rect 231 28328 1607 28362
rect 231 28232 1607 28266
rect 231 28136 1607 28170
rect 231 28040 1607 28074
rect 231 27944 1607 27978
rect 231 27848 1607 27882
rect 231 27752 1607 27786
rect 231 27656 1607 27690
rect 231 27560 1607 27594
rect 231 27464 1607 27498
rect 231 27368 1607 27402
rect 231 27272 1607 27306
rect 231 27176 1607 27210
rect 231 27080 1607 27114
rect 231 26984 1607 27018
rect 231 26888 1607 26922
rect 231 26792 1607 26826
rect 231 26696 1607 26730
rect 231 26600 1607 26634
rect 231 26504 1607 26538
rect 231 26408 1607 26442
rect 231 26312 1607 26346
rect 231 26216 1607 26250
rect 231 26120 1607 26154
rect 231 26024 1607 26058
rect 231 25928 1607 25962
rect 231 25832 1607 25866
rect 231 25736 1607 25770
rect 231 25640 1607 25674
rect 231 25544 1607 25578
rect 231 25448 1607 25482
rect 231 25352 1607 25386
rect 231 25256 1607 25290
rect 231 25160 1607 25194
rect 231 25064 1607 25098
rect 231 24968 1607 25002
rect 231 24872 1607 24906
rect 231 24776 1607 24810
rect 231 24680 1607 24714
rect 231 24584 1607 24618
rect 231 24488 1607 24522
rect 231 24392 1607 24426
rect 231 24296 1607 24330
rect 231 24200 1607 24234
rect 231 24104 1607 24138
rect 231 24008 1607 24042
rect 231 23912 1607 23946
rect 231 23816 1607 23850
rect 231 23720 1607 23754
rect 231 23624 1607 23658
rect 231 23528 1607 23562
rect 231 23432 1607 23466
rect 231 23336 1607 23370
rect 231 23240 1607 23274
rect 231 23144 1607 23178
rect 231 23048 1607 23082
rect 231 21670 1607 21704
rect 231 21574 1607 21608
rect 231 21478 1607 21512
rect 231 21382 1607 21416
rect 231 21286 1607 21320
rect 231 21190 1607 21224
rect 231 21094 1607 21128
rect 231 20998 1607 21032
rect 231 20902 1607 20936
rect 231 20806 1607 20840
rect 231 20710 1607 20744
rect 231 20614 1607 20648
rect 231 20518 1607 20552
rect 231 20422 1607 20456
rect 231 20326 1607 20360
rect 231 20230 1607 20264
rect 231 20134 1607 20168
rect 231 20038 1607 20072
rect 231 19942 1607 19976
rect 231 19846 1607 19880
rect 231 19750 1607 19784
rect 231 19654 1607 19688
rect 231 19558 1607 19592
rect 231 19462 1607 19496
rect 231 19366 1607 19400
rect 231 19270 1607 19304
rect 231 19174 1607 19208
rect 231 19078 1607 19112
rect 231 18982 1607 19016
rect 231 18886 1607 18920
rect 231 18790 1607 18824
rect 231 18694 1607 18728
rect 231 18598 1607 18632
rect 231 18502 1607 18536
rect 231 18406 1607 18440
rect 231 18310 1607 18344
rect 231 18214 1607 18248
rect 231 18118 1607 18152
rect 231 18022 1607 18056
rect 231 17926 1607 17960
rect 231 17830 1607 17864
rect 231 17734 1607 17768
rect 231 17638 1607 17672
rect 231 17542 1607 17576
rect 231 17446 1607 17480
rect 231 17350 1607 17384
rect 231 17254 1607 17288
rect 231 17158 1607 17192
rect 231 17062 1607 17096
rect 231 16966 1607 17000
rect 231 16870 1607 16904
rect 231 16774 1607 16808
rect 231 16678 1607 16712
rect 231 16582 1607 16616
rect 231 16486 1607 16520
rect 231 16390 1607 16424
rect 231 16294 1607 16328
rect 231 16198 1607 16232
rect 231 16102 1607 16136
rect 231 16006 1607 16040
rect 231 15910 1607 15944
rect 231 15814 1607 15848
rect 231 15718 1607 15752
rect 231 15622 1607 15656
rect 231 15526 1607 15560
rect 231 15430 1607 15464
rect 231 15334 1607 15368
rect 231 15238 1607 15272
rect 231 15142 1607 15176
rect 231 15046 1607 15080
rect 231 14950 1607 14984
rect 231 14854 1607 14888
rect 231 14758 1607 14792
rect 231 14662 1607 14696
rect 231 14566 1607 14600
rect 231 14470 1607 14504
rect 231 14374 1607 14408
rect 231 14278 1607 14312
rect 231 14182 1607 14216
rect 231 14086 1607 14120
rect 231 13990 1607 14024
rect 231 13894 1607 13928
rect 231 13798 1607 13832
rect 231 13702 1607 13736
rect 231 13606 1607 13640
rect 231 13510 1607 13544
rect 231 13414 1607 13448
rect 231 13318 1607 13352
rect 231 13222 1607 13256
rect 231 13126 1607 13160
rect 231 13030 1607 13064
rect 231 12934 1607 12968
rect 231 12838 1607 12872
rect 231 12742 1607 12776
rect 231 12646 1607 12680
rect 231 12550 1607 12584
rect 231 12454 1607 12488
rect 231 12358 1607 12392
rect 231 12262 1607 12296
rect 231 12166 1607 12200
rect 231 12070 1607 12104
rect 231 11974 1607 12008
rect 231 11878 1607 11912
rect 231 11782 1607 11816
rect 231 11686 1607 11720
rect 231 11590 1607 11624
rect 231 11494 1607 11528
rect 231 11398 1607 11432
rect 231 11302 1607 11336
rect 231 11206 1607 11240
rect 231 11110 1607 11144
rect 231 11014 1607 11048
rect 231 10918 1607 10952
rect 231 10822 1607 10856
rect 231 10726 1607 10760
rect 231 10630 1607 10664
rect 231 10534 1607 10568
rect 231 10438 1607 10472
rect 231 10342 1607 10376
rect 231 10246 1607 10280
rect 231 10150 1607 10184
rect 231 10054 1607 10088
rect 231 9958 1607 9992
rect 231 9862 1607 9896
rect 231 9766 1607 9800
rect 231 9670 1607 9704
rect 231 9574 1607 9608
rect 231 9478 1607 9512
rect 231 9382 1607 9416
rect 231 9286 1607 9320
rect 231 9190 1607 9224
rect 231 9094 1607 9128
rect 231 8998 1607 9032
rect 231 8902 1607 8936
rect 231 8806 1607 8840
rect 231 8710 1607 8744
rect 231 8614 1607 8648
rect 231 8518 1607 8552
rect 231 8422 1607 8456
rect 231 8326 1607 8360
rect 231 8230 1607 8264
rect 231 8134 1607 8168
rect 231 8038 1607 8072
rect 231 7942 1607 7976
rect 231 7846 1607 7880
rect 231 7750 1607 7784
rect 231 7654 1607 7688
rect 231 7558 1607 7592
rect 231 7462 1607 7496
rect 231 7366 1607 7400
rect 231 7270 1607 7304
rect 231 7174 1607 7208
rect 231 7078 1607 7112
rect 231 6982 1607 7016
rect 231 6886 1607 6920
rect 231 6790 1607 6824
rect 231 6694 1607 6728
rect 231 6598 1607 6632
rect 231 6502 1607 6536
rect 231 6406 1607 6440
rect 231 6310 1607 6344
rect 231 6214 1607 6248
rect 231 6118 1607 6152
rect 231 6022 1607 6056
rect 231 5926 1607 5960
rect 231 5830 1607 5864
rect 231 5734 1607 5768
rect 231 5638 1607 5672
rect 231 5542 1607 5576
rect 231 5446 1607 5480
rect 231 5350 1607 5384
rect 231 5254 1607 5288
rect 231 5158 1607 5192
rect 231 5062 1607 5096
rect 231 4966 1607 5000
rect 231 4870 1607 4904
rect 231 4774 1607 4808
rect 231 4678 1607 4712
rect 231 4582 1607 4616
rect 231 4486 1607 4520
rect 231 4390 1607 4424
rect 231 4294 1607 4328
rect 231 4198 1607 4232
rect 231 4102 1607 4136
rect 231 4006 1607 4040
rect 231 3910 1607 3944
rect 231 3814 1607 3848
rect 231 3718 1607 3752
rect 231 3622 1607 3656
rect 231 3526 1607 3560
rect 231 3430 1607 3464
rect 231 3334 1607 3368
rect 231 3238 1607 3272
rect 231 3142 1607 3176
rect 231 3046 1607 3080
rect 231 2950 1607 2984
rect 231 2854 1607 2888
rect 231 2758 1607 2792
rect 231 2662 1607 2696
rect 231 2566 1607 2600
rect 231 2470 1607 2504
rect 231 2374 1607 2408
rect 231 2278 1607 2312
rect 231 2182 1607 2216
rect 231 2086 1607 2120
rect 231 1990 1607 2024
rect 231 1894 1607 1928
rect 231 1798 1607 1832
rect 231 1702 1607 1736
rect 231 1606 1607 1640
rect 231 1510 1607 1544
rect 231 1414 1607 1448
rect 231 1318 1607 1352
rect 231 1222 1607 1256
rect 231 1126 1607 1160
rect 231 1030 1607 1064
rect 231 934 1607 968
rect 231 838 1607 872
rect 231 742 1607 776
rect 231 646 1607 680
rect 231 550 1607 584
<< nsubdiff >>
rect 36 44282 132 44316
rect 1706 44282 1802 44316
rect 36 44220 70 44282
rect 1768 44220 1802 44282
rect 36 22968 70 23030
rect 1768 22968 1802 23030
rect 36 22934 132 22968
rect 1706 22934 1802 22968
rect 36 21784 132 21818
rect 1706 21784 1802 21818
rect 36 21722 70 21784
rect 1768 21722 1802 21784
rect 36 470 70 532
rect 1768 470 1802 532
rect 36 436 132 470
rect 1706 436 1802 470
<< nsubdiffcont >>
rect 132 44282 1706 44316
rect 36 23030 70 44220
rect 1768 23030 1802 44220
rect 132 22934 1706 22968
rect 132 21784 1706 21818
rect 36 532 70 21722
rect 1768 532 1802 21722
rect 132 436 1706 470
<< poly >>
rect 122 44154 188 44170
rect 122 44120 138 44154
rect 172 44152 188 44154
rect 172 44122 219 44152
rect 1619 44122 1645 44152
rect 172 44120 188 44122
rect 122 44104 188 44120
rect 1650 44058 1716 44074
rect 1650 44056 1666 44058
rect 193 44026 219 44056
rect 1619 44026 1666 44056
rect 122 43962 188 43978
rect 122 43928 138 43962
rect 172 43960 188 43962
rect 1650 44024 1666 44026
rect 1700 44024 1716 44058
rect 1650 44008 1716 44024
rect 172 43930 219 43960
rect 1619 43930 1645 43960
rect 172 43928 188 43930
rect 122 43912 188 43928
rect 1650 43866 1716 43882
rect 1650 43864 1666 43866
rect 193 43834 219 43864
rect 1619 43834 1666 43864
rect 122 43770 188 43786
rect 122 43736 138 43770
rect 172 43768 188 43770
rect 1650 43832 1666 43834
rect 1700 43832 1716 43866
rect 1650 43816 1716 43832
rect 172 43738 219 43768
rect 1619 43738 1645 43768
rect 172 43736 188 43738
rect 122 43720 188 43736
rect 1650 43674 1716 43690
rect 1650 43672 1666 43674
rect 193 43642 219 43672
rect 1619 43642 1666 43672
rect 122 43578 188 43594
rect 122 43544 138 43578
rect 172 43576 188 43578
rect 1650 43640 1666 43642
rect 1700 43640 1716 43674
rect 1650 43624 1716 43640
rect 172 43546 219 43576
rect 1619 43546 1645 43576
rect 172 43544 188 43546
rect 122 43528 188 43544
rect 1650 43482 1716 43498
rect 1650 43480 1666 43482
rect 193 43450 219 43480
rect 1619 43450 1666 43480
rect 122 43386 188 43402
rect 122 43352 138 43386
rect 172 43384 188 43386
rect 1650 43448 1666 43450
rect 1700 43448 1716 43482
rect 1650 43432 1716 43448
rect 172 43354 219 43384
rect 1619 43354 1645 43384
rect 172 43352 188 43354
rect 122 43336 188 43352
rect 1650 43290 1716 43306
rect 1650 43288 1666 43290
rect 193 43258 219 43288
rect 1619 43258 1666 43288
rect 122 43194 188 43210
rect 122 43160 138 43194
rect 172 43192 188 43194
rect 1650 43256 1666 43258
rect 1700 43256 1716 43290
rect 1650 43240 1716 43256
rect 172 43162 219 43192
rect 1619 43162 1645 43192
rect 172 43160 188 43162
rect 122 43144 188 43160
rect 1650 43098 1716 43114
rect 1650 43096 1666 43098
rect 193 43066 219 43096
rect 1619 43066 1666 43096
rect 122 43002 188 43018
rect 122 42968 138 43002
rect 172 43000 188 43002
rect 1650 43064 1666 43066
rect 1700 43064 1716 43098
rect 1650 43048 1716 43064
rect 172 42970 219 43000
rect 1619 42970 1645 43000
rect 172 42968 188 42970
rect 122 42952 188 42968
rect 1650 42906 1716 42922
rect 1650 42904 1666 42906
rect 193 42874 219 42904
rect 1619 42874 1666 42904
rect 122 42810 188 42826
rect 122 42776 138 42810
rect 172 42808 188 42810
rect 1650 42872 1666 42874
rect 1700 42872 1716 42906
rect 1650 42856 1716 42872
rect 172 42778 219 42808
rect 1619 42778 1645 42808
rect 172 42776 188 42778
rect 122 42760 188 42776
rect 1650 42714 1716 42730
rect 1650 42712 1666 42714
rect 193 42682 219 42712
rect 1619 42682 1666 42712
rect 122 42618 188 42634
rect 122 42584 138 42618
rect 172 42616 188 42618
rect 1650 42680 1666 42682
rect 1700 42680 1716 42714
rect 1650 42664 1716 42680
rect 172 42586 219 42616
rect 1619 42586 1645 42616
rect 172 42584 188 42586
rect 122 42568 188 42584
rect 1650 42522 1716 42538
rect 1650 42520 1666 42522
rect 193 42490 219 42520
rect 1619 42490 1666 42520
rect 122 42426 188 42442
rect 122 42392 138 42426
rect 172 42424 188 42426
rect 1650 42488 1666 42490
rect 1700 42488 1716 42522
rect 1650 42472 1716 42488
rect 172 42394 219 42424
rect 1619 42394 1645 42424
rect 172 42392 188 42394
rect 122 42376 188 42392
rect 1650 42330 1716 42346
rect 1650 42328 1666 42330
rect 193 42298 219 42328
rect 1619 42298 1666 42328
rect 122 42234 188 42250
rect 122 42200 138 42234
rect 172 42232 188 42234
rect 1650 42296 1666 42298
rect 1700 42296 1716 42330
rect 1650 42280 1716 42296
rect 172 42202 219 42232
rect 1619 42202 1645 42232
rect 172 42200 188 42202
rect 122 42184 188 42200
rect 1650 42138 1716 42154
rect 1650 42136 1666 42138
rect 193 42106 219 42136
rect 1619 42106 1666 42136
rect 122 42042 188 42058
rect 122 42008 138 42042
rect 172 42040 188 42042
rect 1650 42104 1666 42106
rect 1700 42104 1716 42138
rect 1650 42088 1716 42104
rect 172 42010 219 42040
rect 1619 42010 1645 42040
rect 172 42008 188 42010
rect 122 41992 188 42008
rect 1650 41946 1716 41962
rect 1650 41944 1666 41946
rect 193 41914 219 41944
rect 1619 41914 1666 41944
rect 122 41850 188 41866
rect 122 41816 138 41850
rect 172 41848 188 41850
rect 1650 41912 1666 41914
rect 1700 41912 1716 41946
rect 1650 41896 1716 41912
rect 172 41818 219 41848
rect 1619 41818 1645 41848
rect 172 41816 188 41818
rect 122 41800 188 41816
rect 1650 41754 1716 41770
rect 1650 41752 1666 41754
rect 193 41722 219 41752
rect 1619 41722 1666 41752
rect 122 41658 188 41674
rect 122 41624 138 41658
rect 172 41656 188 41658
rect 1650 41720 1666 41722
rect 1700 41720 1716 41754
rect 1650 41704 1716 41720
rect 172 41626 219 41656
rect 1619 41626 1645 41656
rect 172 41624 188 41626
rect 122 41608 188 41624
rect 1650 41562 1716 41578
rect 1650 41560 1666 41562
rect 193 41530 219 41560
rect 1619 41530 1666 41560
rect 122 41466 188 41482
rect 122 41432 138 41466
rect 172 41464 188 41466
rect 1650 41528 1666 41530
rect 1700 41528 1716 41562
rect 1650 41512 1716 41528
rect 172 41434 219 41464
rect 1619 41434 1645 41464
rect 172 41432 188 41434
rect 122 41416 188 41432
rect 1650 41370 1716 41386
rect 1650 41368 1666 41370
rect 193 41338 219 41368
rect 1619 41338 1666 41368
rect 122 41274 188 41290
rect 122 41240 138 41274
rect 172 41272 188 41274
rect 1650 41336 1666 41338
rect 1700 41336 1716 41370
rect 1650 41320 1716 41336
rect 172 41242 219 41272
rect 1619 41242 1645 41272
rect 172 41240 188 41242
rect 122 41224 188 41240
rect 1650 41178 1716 41194
rect 1650 41176 1666 41178
rect 193 41146 219 41176
rect 1619 41146 1666 41176
rect 122 41082 188 41098
rect 122 41048 138 41082
rect 172 41080 188 41082
rect 1650 41144 1666 41146
rect 1700 41144 1716 41178
rect 1650 41128 1716 41144
rect 172 41050 219 41080
rect 1619 41050 1645 41080
rect 172 41048 188 41050
rect 122 41032 188 41048
rect 1650 40986 1716 41002
rect 1650 40984 1666 40986
rect 193 40954 219 40984
rect 1619 40954 1666 40984
rect 122 40890 188 40906
rect 122 40856 138 40890
rect 172 40888 188 40890
rect 1650 40952 1666 40954
rect 1700 40952 1716 40986
rect 1650 40936 1716 40952
rect 172 40858 219 40888
rect 1619 40858 1645 40888
rect 172 40856 188 40858
rect 122 40840 188 40856
rect 1650 40794 1716 40810
rect 1650 40792 1666 40794
rect 193 40762 219 40792
rect 1619 40762 1666 40792
rect 122 40698 188 40714
rect 122 40664 138 40698
rect 172 40696 188 40698
rect 1650 40760 1666 40762
rect 1700 40760 1716 40794
rect 1650 40744 1716 40760
rect 172 40666 219 40696
rect 1619 40666 1645 40696
rect 172 40664 188 40666
rect 122 40648 188 40664
rect 1650 40602 1716 40618
rect 1650 40600 1666 40602
rect 193 40570 219 40600
rect 1619 40570 1666 40600
rect 122 40506 188 40522
rect 122 40472 138 40506
rect 172 40504 188 40506
rect 1650 40568 1666 40570
rect 1700 40568 1716 40602
rect 1650 40552 1716 40568
rect 172 40474 219 40504
rect 1619 40474 1645 40504
rect 172 40472 188 40474
rect 122 40456 188 40472
rect 1650 40410 1716 40426
rect 1650 40408 1666 40410
rect 193 40378 219 40408
rect 1619 40378 1666 40408
rect 122 40314 188 40330
rect 122 40280 138 40314
rect 172 40312 188 40314
rect 1650 40376 1666 40378
rect 1700 40376 1716 40410
rect 1650 40360 1716 40376
rect 172 40282 219 40312
rect 1619 40282 1645 40312
rect 172 40280 188 40282
rect 122 40264 188 40280
rect 1650 40218 1716 40234
rect 1650 40216 1666 40218
rect 193 40186 219 40216
rect 1619 40186 1666 40216
rect 122 40122 188 40138
rect 122 40088 138 40122
rect 172 40120 188 40122
rect 1650 40184 1666 40186
rect 1700 40184 1716 40218
rect 1650 40168 1716 40184
rect 172 40090 219 40120
rect 1619 40090 1645 40120
rect 172 40088 188 40090
rect 122 40072 188 40088
rect 1650 40026 1716 40042
rect 1650 40024 1666 40026
rect 193 39994 219 40024
rect 1619 39994 1666 40024
rect 122 39930 188 39946
rect 122 39896 138 39930
rect 172 39928 188 39930
rect 1650 39992 1666 39994
rect 1700 39992 1716 40026
rect 1650 39976 1716 39992
rect 172 39898 219 39928
rect 1619 39898 1645 39928
rect 172 39896 188 39898
rect 122 39880 188 39896
rect 1650 39834 1716 39850
rect 1650 39832 1666 39834
rect 193 39802 219 39832
rect 1619 39802 1666 39832
rect 122 39738 188 39754
rect 122 39704 138 39738
rect 172 39736 188 39738
rect 1650 39800 1666 39802
rect 1700 39800 1716 39834
rect 1650 39784 1716 39800
rect 172 39706 219 39736
rect 1619 39706 1645 39736
rect 172 39704 188 39706
rect 122 39688 188 39704
rect 1650 39642 1716 39658
rect 1650 39640 1666 39642
rect 193 39610 219 39640
rect 1619 39610 1666 39640
rect 122 39546 188 39562
rect 122 39512 138 39546
rect 172 39544 188 39546
rect 1650 39608 1666 39610
rect 1700 39608 1716 39642
rect 1650 39592 1716 39608
rect 172 39514 219 39544
rect 1619 39514 1645 39544
rect 172 39512 188 39514
rect 122 39496 188 39512
rect 1650 39450 1716 39466
rect 1650 39448 1666 39450
rect 193 39418 219 39448
rect 1619 39418 1666 39448
rect 122 39354 188 39370
rect 122 39320 138 39354
rect 172 39352 188 39354
rect 1650 39416 1666 39418
rect 1700 39416 1716 39450
rect 1650 39400 1716 39416
rect 172 39322 219 39352
rect 1619 39322 1645 39352
rect 172 39320 188 39322
rect 122 39304 188 39320
rect 1650 39258 1716 39274
rect 1650 39256 1666 39258
rect 193 39226 219 39256
rect 1619 39226 1666 39256
rect 122 39162 188 39178
rect 122 39128 138 39162
rect 172 39160 188 39162
rect 1650 39224 1666 39226
rect 1700 39224 1716 39258
rect 1650 39208 1716 39224
rect 172 39130 219 39160
rect 1619 39130 1645 39160
rect 172 39128 188 39130
rect 122 39112 188 39128
rect 1650 39066 1716 39082
rect 1650 39064 1666 39066
rect 193 39034 219 39064
rect 1619 39034 1666 39064
rect 122 38970 188 38986
rect 122 38936 138 38970
rect 172 38968 188 38970
rect 1650 39032 1666 39034
rect 1700 39032 1716 39066
rect 1650 39016 1716 39032
rect 172 38938 219 38968
rect 1619 38938 1645 38968
rect 172 38936 188 38938
rect 122 38920 188 38936
rect 1650 38874 1716 38890
rect 1650 38872 1666 38874
rect 193 38842 219 38872
rect 1619 38842 1666 38872
rect 122 38778 188 38794
rect 122 38744 138 38778
rect 172 38776 188 38778
rect 1650 38840 1666 38842
rect 1700 38840 1716 38874
rect 1650 38824 1716 38840
rect 172 38746 219 38776
rect 1619 38746 1645 38776
rect 172 38744 188 38746
rect 122 38728 188 38744
rect 1650 38682 1716 38698
rect 1650 38680 1666 38682
rect 193 38650 219 38680
rect 1619 38650 1666 38680
rect 122 38586 188 38602
rect 122 38552 138 38586
rect 172 38584 188 38586
rect 1650 38648 1666 38650
rect 1700 38648 1716 38682
rect 1650 38632 1716 38648
rect 172 38554 219 38584
rect 1619 38554 1645 38584
rect 172 38552 188 38554
rect 122 38536 188 38552
rect 1650 38490 1716 38506
rect 1650 38488 1666 38490
rect 193 38458 219 38488
rect 1619 38458 1666 38488
rect 122 38394 188 38410
rect 122 38360 138 38394
rect 172 38392 188 38394
rect 1650 38456 1666 38458
rect 1700 38456 1716 38490
rect 1650 38440 1716 38456
rect 172 38362 219 38392
rect 1619 38362 1645 38392
rect 172 38360 188 38362
rect 122 38344 188 38360
rect 1650 38298 1716 38314
rect 1650 38296 1666 38298
rect 193 38266 219 38296
rect 1619 38266 1666 38296
rect 122 38202 188 38218
rect 122 38168 138 38202
rect 172 38200 188 38202
rect 1650 38264 1666 38266
rect 1700 38264 1716 38298
rect 1650 38248 1716 38264
rect 172 38170 219 38200
rect 1619 38170 1645 38200
rect 172 38168 188 38170
rect 122 38152 188 38168
rect 1650 38106 1716 38122
rect 1650 38104 1666 38106
rect 193 38074 219 38104
rect 1619 38074 1666 38104
rect 122 38010 188 38026
rect 122 37976 138 38010
rect 172 38008 188 38010
rect 1650 38072 1666 38074
rect 1700 38072 1716 38106
rect 1650 38056 1716 38072
rect 172 37978 219 38008
rect 1619 37978 1645 38008
rect 172 37976 188 37978
rect 122 37960 188 37976
rect 1650 37914 1716 37930
rect 1650 37912 1666 37914
rect 193 37882 219 37912
rect 1619 37882 1666 37912
rect 122 37818 188 37834
rect 122 37784 138 37818
rect 172 37816 188 37818
rect 1650 37880 1666 37882
rect 1700 37880 1716 37914
rect 1650 37864 1716 37880
rect 172 37786 219 37816
rect 1619 37786 1645 37816
rect 172 37784 188 37786
rect 122 37768 188 37784
rect 1650 37722 1716 37738
rect 1650 37720 1666 37722
rect 193 37690 219 37720
rect 1619 37690 1666 37720
rect 122 37626 188 37642
rect 122 37592 138 37626
rect 172 37624 188 37626
rect 1650 37688 1666 37690
rect 1700 37688 1716 37722
rect 1650 37672 1716 37688
rect 172 37594 219 37624
rect 1619 37594 1645 37624
rect 172 37592 188 37594
rect 122 37576 188 37592
rect 1650 37530 1716 37546
rect 1650 37528 1666 37530
rect 193 37498 219 37528
rect 1619 37498 1666 37528
rect 122 37434 188 37450
rect 122 37400 138 37434
rect 172 37432 188 37434
rect 1650 37496 1666 37498
rect 1700 37496 1716 37530
rect 1650 37480 1716 37496
rect 172 37402 219 37432
rect 1619 37402 1645 37432
rect 172 37400 188 37402
rect 122 37384 188 37400
rect 1650 37338 1716 37354
rect 1650 37336 1666 37338
rect 193 37306 219 37336
rect 1619 37306 1666 37336
rect 122 37242 188 37258
rect 122 37208 138 37242
rect 172 37240 188 37242
rect 1650 37304 1666 37306
rect 1700 37304 1716 37338
rect 1650 37288 1716 37304
rect 172 37210 219 37240
rect 1619 37210 1645 37240
rect 172 37208 188 37210
rect 122 37192 188 37208
rect 1650 37146 1716 37162
rect 1650 37144 1666 37146
rect 193 37114 219 37144
rect 1619 37114 1666 37144
rect 122 37050 188 37066
rect 122 37016 138 37050
rect 172 37048 188 37050
rect 1650 37112 1666 37114
rect 1700 37112 1716 37146
rect 1650 37096 1716 37112
rect 172 37018 219 37048
rect 1619 37018 1645 37048
rect 172 37016 188 37018
rect 122 37000 188 37016
rect 1650 36954 1716 36970
rect 1650 36952 1666 36954
rect 193 36922 219 36952
rect 1619 36922 1666 36952
rect 122 36858 188 36874
rect 122 36824 138 36858
rect 172 36856 188 36858
rect 1650 36920 1666 36922
rect 1700 36920 1716 36954
rect 1650 36904 1716 36920
rect 172 36826 219 36856
rect 1619 36826 1645 36856
rect 172 36824 188 36826
rect 122 36808 188 36824
rect 1650 36762 1716 36778
rect 1650 36760 1666 36762
rect 193 36730 219 36760
rect 1619 36730 1666 36760
rect 122 36666 188 36682
rect 122 36632 138 36666
rect 172 36664 188 36666
rect 1650 36728 1666 36730
rect 1700 36728 1716 36762
rect 1650 36712 1716 36728
rect 172 36634 219 36664
rect 1619 36634 1645 36664
rect 172 36632 188 36634
rect 122 36616 188 36632
rect 1650 36570 1716 36586
rect 1650 36568 1666 36570
rect 193 36538 219 36568
rect 1619 36538 1666 36568
rect 122 36474 188 36490
rect 122 36440 138 36474
rect 172 36472 188 36474
rect 1650 36536 1666 36538
rect 1700 36536 1716 36570
rect 1650 36520 1716 36536
rect 172 36442 219 36472
rect 1619 36442 1645 36472
rect 172 36440 188 36442
rect 122 36424 188 36440
rect 1650 36378 1716 36394
rect 1650 36376 1666 36378
rect 193 36346 219 36376
rect 1619 36346 1666 36376
rect 122 36282 188 36298
rect 122 36248 138 36282
rect 172 36280 188 36282
rect 1650 36344 1666 36346
rect 1700 36344 1716 36378
rect 1650 36328 1716 36344
rect 172 36250 219 36280
rect 1619 36250 1645 36280
rect 172 36248 188 36250
rect 122 36232 188 36248
rect 1650 36186 1716 36202
rect 1650 36184 1666 36186
rect 193 36154 219 36184
rect 1619 36154 1666 36184
rect 122 36090 188 36106
rect 122 36056 138 36090
rect 172 36088 188 36090
rect 1650 36152 1666 36154
rect 1700 36152 1716 36186
rect 1650 36136 1716 36152
rect 172 36058 219 36088
rect 1619 36058 1645 36088
rect 172 36056 188 36058
rect 122 36040 188 36056
rect 1650 35994 1716 36010
rect 1650 35992 1666 35994
rect 193 35962 219 35992
rect 1619 35962 1666 35992
rect 122 35898 188 35914
rect 122 35864 138 35898
rect 172 35896 188 35898
rect 1650 35960 1666 35962
rect 1700 35960 1716 35994
rect 1650 35944 1716 35960
rect 172 35866 219 35896
rect 1619 35866 1645 35896
rect 172 35864 188 35866
rect 122 35848 188 35864
rect 1650 35802 1716 35818
rect 1650 35800 1666 35802
rect 193 35770 219 35800
rect 1619 35770 1666 35800
rect 122 35706 188 35722
rect 122 35672 138 35706
rect 172 35704 188 35706
rect 1650 35768 1666 35770
rect 1700 35768 1716 35802
rect 1650 35752 1716 35768
rect 172 35674 219 35704
rect 1619 35674 1645 35704
rect 172 35672 188 35674
rect 122 35656 188 35672
rect 1650 35610 1716 35626
rect 1650 35608 1666 35610
rect 193 35578 219 35608
rect 1619 35578 1666 35608
rect 122 35514 188 35530
rect 122 35480 138 35514
rect 172 35512 188 35514
rect 1650 35576 1666 35578
rect 1700 35576 1716 35610
rect 1650 35560 1716 35576
rect 172 35482 219 35512
rect 1619 35482 1645 35512
rect 172 35480 188 35482
rect 122 35464 188 35480
rect 1650 35418 1716 35434
rect 1650 35416 1666 35418
rect 193 35386 219 35416
rect 1619 35386 1666 35416
rect 122 35322 188 35338
rect 122 35288 138 35322
rect 172 35320 188 35322
rect 1650 35384 1666 35386
rect 1700 35384 1716 35418
rect 1650 35368 1716 35384
rect 172 35290 219 35320
rect 1619 35290 1645 35320
rect 172 35288 188 35290
rect 122 35272 188 35288
rect 1650 35226 1716 35242
rect 1650 35224 1666 35226
rect 193 35194 219 35224
rect 1619 35194 1666 35224
rect 122 35130 188 35146
rect 122 35096 138 35130
rect 172 35128 188 35130
rect 1650 35192 1666 35194
rect 1700 35192 1716 35226
rect 1650 35176 1716 35192
rect 172 35098 219 35128
rect 1619 35098 1645 35128
rect 172 35096 188 35098
rect 122 35080 188 35096
rect 1650 35034 1716 35050
rect 1650 35032 1666 35034
rect 193 35002 219 35032
rect 1619 35002 1666 35032
rect 122 34938 188 34954
rect 122 34904 138 34938
rect 172 34936 188 34938
rect 1650 35000 1666 35002
rect 1700 35000 1716 35034
rect 1650 34984 1716 35000
rect 172 34906 219 34936
rect 1619 34906 1645 34936
rect 172 34904 188 34906
rect 122 34888 188 34904
rect 1650 34842 1716 34858
rect 1650 34840 1666 34842
rect 193 34810 219 34840
rect 1619 34810 1666 34840
rect 122 34746 188 34762
rect 122 34712 138 34746
rect 172 34744 188 34746
rect 1650 34808 1666 34810
rect 1700 34808 1716 34842
rect 1650 34792 1716 34808
rect 172 34714 219 34744
rect 1619 34714 1645 34744
rect 172 34712 188 34714
rect 122 34696 188 34712
rect 1650 34650 1716 34666
rect 1650 34648 1666 34650
rect 193 34618 219 34648
rect 1619 34618 1666 34648
rect 122 34554 188 34570
rect 122 34520 138 34554
rect 172 34552 188 34554
rect 1650 34616 1666 34618
rect 1700 34616 1716 34650
rect 1650 34600 1716 34616
rect 172 34522 219 34552
rect 1619 34522 1645 34552
rect 172 34520 188 34522
rect 122 34504 188 34520
rect 1650 34458 1716 34474
rect 1650 34456 1666 34458
rect 193 34426 219 34456
rect 1619 34426 1666 34456
rect 122 34362 188 34378
rect 122 34328 138 34362
rect 172 34360 188 34362
rect 1650 34424 1666 34426
rect 1700 34424 1716 34458
rect 1650 34408 1716 34424
rect 172 34330 219 34360
rect 1619 34330 1645 34360
rect 172 34328 188 34330
rect 122 34312 188 34328
rect 1650 34266 1716 34282
rect 1650 34264 1666 34266
rect 193 34234 219 34264
rect 1619 34234 1666 34264
rect 122 34170 188 34186
rect 122 34136 138 34170
rect 172 34168 188 34170
rect 1650 34232 1666 34234
rect 1700 34232 1716 34266
rect 1650 34216 1716 34232
rect 172 34138 219 34168
rect 1619 34138 1645 34168
rect 172 34136 188 34138
rect 122 34120 188 34136
rect 1650 34074 1716 34090
rect 1650 34072 1666 34074
rect 193 34042 219 34072
rect 1619 34042 1666 34072
rect 122 33978 188 33994
rect 122 33944 138 33978
rect 172 33976 188 33978
rect 1650 34040 1666 34042
rect 1700 34040 1716 34074
rect 1650 34024 1716 34040
rect 172 33946 219 33976
rect 1619 33946 1645 33976
rect 172 33944 188 33946
rect 122 33928 188 33944
rect 1650 33882 1716 33898
rect 1650 33880 1666 33882
rect 193 33850 219 33880
rect 1619 33850 1666 33880
rect 122 33786 188 33802
rect 122 33752 138 33786
rect 172 33784 188 33786
rect 1650 33848 1666 33850
rect 1700 33848 1716 33882
rect 1650 33832 1716 33848
rect 172 33754 219 33784
rect 1619 33754 1645 33784
rect 172 33752 188 33754
rect 122 33736 188 33752
rect 1650 33690 1716 33706
rect 1650 33688 1666 33690
rect 193 33658 219 33688
rect 1619 33658 1666 33688
rect 122 33594 188 33610
rect 122 33560 138 33594
rect 172 33592 188 33594
rect 1650 33656 1666 33658
rect 1700 33656 1716 33690
rect 1650 33640 1716 33656
rect 172 33562 219 33592
rect 1619 33562 1645 33592
rect 172 33560 188 33562
rect 122 33544 188 33560
rect 1650 33498 1716 33514
rect 1650 33496 1666 33498
rect 193 33466 219 33496
rect 1619 33466 1666 33496
rect 122 33402 188 33418
rect 122 33368 138 33402
rect 172 33400 188 33402
rect 1650 33464 1666 33466
rect 1700 33464 1716 33498
rect 1650 33448 1716 33464
rect 172 33370 219 33400
rect 1619 33370 1645 33400
rect 172 33368 188 33370
rect 122 33352 188 33368
rect 1650 33306 1716 33322
rect 1650 33304 1666 33306
rect 193 33274 219 33304
rect 1619 33274 1666 33304
rect 122 33210 188 33226
rect 122 33176 138 33210
rect 172 33208 188 33210
rect 1650 33272 1666 33274
rect 1700 33272 1716 33306
rect 1650 33256 1716 33272
rect 172 33178 219 33208
rect 1619 33178 1645 33208
rect 172 33176 188 33178
rect 122 33160 188 33176
rect 1650 33114 1716 33130
rect 1650 33112 1666 33114
rect 193 33082 219 33112
rect 1619 33082 1666 33112
rect 122 33018 188 33034
rect 122 32984 138 33018
rect 172 33016 188 33018
rect 1650 33080 1666 33082
rect 1700 33080 1716 33114
rect 1650 33064 1716 33080
rect 172 32986 219 33016
rect 1619 32986 1645 33016
rect 172 32984 188 32986
rect 122 32968 188 32984
rect 1650 32922 1716 32938
rect 1650 32920 1666 32922
rect 193 32890 219 32920
rect 1619 32890 1666 32920
rect 122 32826 188 32842
rect 122 32792 138 32826
rect 172 32824 188 32826
rect 1650 32888 1666 32890
rect 1700 32888 1716 32922
rect 1650 32872 1716 32888
rect 172 32794 219 32824
rect 1619 32794 1645 32824
rect 172 32792 188 32794
rect 122 32776 188 32792
rect 1650 32730 1716 32746
rect 1650 32728 1666 32730
rect 193 32698 219 32728
rect 1619 32698 1666 32728
rect 122 32634 188 32650
rect 122 32600 138 32634
rect 172 32632 188 32634
rect 1650 32696 1666 32698
rect 1700 32696 1716 32730
rect 1650 32680 1716 32696
rect 172 32602 219 32632
rect 1619 32602 1645 32632
rect 172 32600 188 32602
rect 122 32584 188 32600
rect 1650 32538 1716 32554
rect 1650 32536 1666 32538
rect 193 32506 219 32536
rect 1619 32506 1666 32536
rect 122 32442 188 32458
rect 122 32408 138 32442
rect 172 32440 188 32442
rect 1650 32504 1666 32506
rect 1700 32504 1716 32538
rect 1650 32488 1716 32504
rect 172 32410 219 32440
rect 1619 32410 1645 32440
rect 172 32408 188 32410
rect 122 32392 188 32408
rect 1650 32346 1716 32362
rect 1650 32344 1666 32346
rect 193 32314 219 32344
rect 1619 32314 1666 32344
rect 122 32250 188 32266
rect 122 32216 138 32250
rect 172 32248 188 32250
rect 1650 32312 1666 32314
rect 1700 32312 1716 32346
rect 1650 32296 1716 32312
rect 172 32218 219 32248
rect 1619 32218 1645 32248
rect 172 32216 188 32218
rect 122 32200 188 32216
rect 1650 32154 1716 32170
rect 1650 32152 1666 32154
rect 193 32122 219 32152
rect 1619 32122 1666 32152
rect 122 32058 188 32074
rect 122 32024 138 32058
rect 172 32056 188 32058
rect 1650 32120 1666 32122
rect 1700 32120 1716 32154
rect 1650 32104 1716 32120
rect 172 32026 219 32056
rect 1619 32026 1645 32056
rect 172 32024 188 32026
rect 122 32008 188 32024
rect 1650 31962 1716 31978
rect 1650 31960 1666 31962
rect 193 31930 219 31960
rect 1619 31930 1666 31960
rect 122 31866 188 31882
rect 122 31832 138 31866
rect 172 31864 188 31866
rect 1650 31928 1666 31930
rect 1700 31928 1716 31962
rect 1650 31912 1716 31928
rect 172 31834 219 31864
rect 1619 31834 1645 31864
rect 172 31832 188 31834
rect 122 31816 188 31832
rect 1650 31770 1716 31786
rect 1650 31768 1666 31770
rect 193 31738 219 31768
rect 1619 31738 1666 31768
rect 122 31674 188 31690
rect 122 31640 138 31674
rect 172 31672 188 31674
rect 1650 31736 1666 31738
rect 1700 31736 1716 31770
rect 1650 31720 1716 31736
rect 172 31642 219 31672
rect 1619 31642 1645 31672
rect 172 31640 188 31642
rect 122 31624 188 31640
rect 1650 31578 1716 31594
rect 1650 31576 1666 31578
rect 193 31546 219 31576
rect 1619 31546 1666 31576
rect 122 31482 188 31498
rect 122 31448 138 31482
rect 172 31480 188 31482
rect 1650 31544 1666 31546
rect 1700 31544 1716 31578
rect 1650 31528 1716 31544
rect 172 31450 219 31480
rect 1619 31450 1645 31480
rect 172 31448 188 31450
rect 122 31432 188 31448
rect 1650 31386 1716 31402
rect 1650 31384 1666 31386
rect 193 31354 219 31384
rect 1619 31354 1666 31384
rect 122 31290 188 31306
rect 122 31256 138 31290
rect 172 31288 188 31290
rect 1650 31352 1666 31354
rect 1700 31352 1716 31386
rect 1650 31336 1716 31352
rect 172 31258 219 31288
rect 1619 31258 1645 31288
rect 172 31256 188 31258
rect 122 31240 188 31256
rect 1650 31194 1716 31210
rect 1650 31192 1666 31194
rect 193 31162 219 31192
rect 1619 31162 1666 31192
rect 122 31098 188 31114
rect 122 31064 138 31098
rect 172 31096 188 31098
rect 1650 31160 1666 31162
rect 1700 31160 1716 31194
rect 1650 31144 1716 31160
rect 172 31066 219 31096
rect 1619 31066 1645 31096
rect 172 31064 188 31066
rect 122 31048 188 31064
rect 1650 31002 1716 31018
rect 1650 31000 1666 31002
rect 193 30970 219 31000
rect 1619 30970 1666 31000
rect 122 30906 188 30922
rect 122 30872 138 30906
rect 172 30904 188 30906
rect 1650 30968 1666 30970
rect 1700 30968 1716 31002
rect 1650 30952 1716 30968
rect 172 30874 219 30904
rect 1619 30874 1645 30904
rect 172 30872 188 30874
rect 122 30856 188 30872
rect 1650 30810 1716 30826
rect 1650 30808 1666 30810
rect 193 30778 219 30808
rect 1619 30778 1666 30808
rect 122 30714 188 30730
rect 122 30680 138 30714
rect 172 30712 188 30714
rect 1650 30776 1666 30778
rect 1700 30776 1716 30810
rect 1650 30760 1716 30776
rect 172 30682 219 30712
rect 1619 30682 1645 30712
rect 172 30680 188 30682
rect 122 30664 188 30680
rect 1650 30618 1716 30634
rect 1650 30616 1666 30618
rect 193 30586 219 30616
rect 1619 30586 1666 30616
rect 122 30522 188 30538
rect 122 30488 138 30522
rect 172 30520 188 30522
rect 1650 30584 1666 30586
rect 1700 30584 1716 30618
rect 1650 30568 1716 30584
rect 172 30490 219 30520
rect 1619 30490 1645 30520
rect 172 30488 188 30490
rect 122 30472 188 30488
rect 1650 30426 1716 30442
rect 1650 30424 1666 30426
rect 193 30394 219 30424
rect 1619 30394 1666 30424
rect 122 30330 188 30346
rect 122 30296 138 30330
rect 172 30328 188 30330
rect 1650 30392 1666 30394
rect 1700 30392 1716 30426
rect 1650 30376 1716 30392
rect 172 30298 219 30328
rect 1619 30298 1645 30328
rect 172 30296 188 30298
rect 122 30280 188 30296
rect 1650 30234 1716 30250
rect 1650 30232 1666 30234
rect 193 30202 219 30232
rect 1619 30202 1666 30232
rect 122 30138 188 30154
rect 122 30104 138 30138
rect 172 30136 188 30138
rect 1650 30200 1666 30202
rect 1700 30200 1716 30234
rect 1650 30184 1716 30200
rect 172 30106 219 30136
rect 1619 30106 1645 30136
rect 172 30104 188 30106
rect 122 30088 188 30104
rect 1650 30042 1716 30058
rect 1650 30040 1666 30042
rect 193 30010 219 30040
rect 1619 30010 1666 30040
rect 122 29946 188 29962
rect 122 29912 138 29946
rect 172 29944 188 29946
rect 1650 30008 1666 30010
rect 1700 30008 1716 30042
rect 1650 29992 1716 30008
rect 172 29914 219 29944
rect 1619 29914 1645 29944
rect 172 29912 188 29914
rect 122 29896 188 29912
rect 1650 29850 1716 29866
rect 1650 29848 1666 29850
rect 193 29818 219 29848
rect 1619 29818 1666 29848
rect 122 29754 188 29770
rect 122 29720 138 29754
rect 172 29752 188 29754
rect 1650 29816 1666 29818
rect 1700 29816 1716 29850
rect 1650 29800 1716 29816
rect 172 29722 219 29752
rect 1619 29722 1645 29752
rect 172 29720 188 29722
rect 122 29704 188 29720
rect 1650 29658 1716 29674
rect 1650 29656 1666 29658
rect 193 29626 219 29656
rect 1619 29626 1666 29656
rect 122 29562 188 29578
rect 122 29528 138 29562
rect 172 29560 188 29562
rect 1650 29624 1666 29626
rect 1700 29624 1716 29658
rect 1650 29608 1716 29624
rect 172 29530 219 29560
rect 1619 29530 1645 29560
rect 172 29528 188 29530
rect 122 29512 188 29528
rect 1650 29466 1716 29482
rect 1650 29464 1666 29466
rect 193 29434 219 29464
rect 1619 29434 1666 29464
rect 122 29370 188 29386
rect 122 29336 138 29370
rect 172 29368 188 29370
rect 1650 29432 1666 29434
rect 1700 29432 1716 29466
rect 1650 29416 1716 29432
rect 172 29338 219 29368
rect 1619 29338 1645 29368
rect 172 29336 188 29338
rect 122 29320 188 29336
rect 1650 29274 1716 29290
rect 1650 29272 1666 29274
rect 193 29242 219 29272
rect 1619 29242 1666 29272
rect 122 29178 188 29194
rect 122 29144 138 29178
rect 172 29176 188 29178
rect 1650 29240 1666 29242
rect 1700 29240 1716 29274
rect 1650 29224 1716 29240
rect 172 29146 219 29176
rect 1619 29146 1645 29176
rect 172 29144 188 29146
rect 122 29128 188 29144
rect 1650 29082 1716 29098
rect 1650 29080 1666 29082
rect 193 29050 219 29080
rect 1619 29050 1666 29080
rect 122 28986 188 29002
rect 122 28952 138 28986
rect 172 28984 188 28986
rect 1650 29048 1666 29050
rect 1700 29048 1716 29082
rect 1650 29032 1716 29048
rect 172 28954 219 28984
rect 1619 28954 1645 28984
rect 172 28952 188 28954
rect 122 28936 188 28952
rect 1650 28890 1716 28906
rect 1650 28888 1666 28890
rect 193 28858 219 28888
rect 1619 28858 1666 28888
rect 122 28794 188 28810
rect 122 28760 138 28794
rect 172 28792 188 28794
rect 1650 28856 1666 28858
rect 1700 28856 1716 28890
rect 1650 28840 1716 28856
rect 172 28762 219 28792
rect 1619 28762 1645 28792
rect 172 28760 188 28762
rect 122 28744 188 28760
rect 1650 28698 1716 28714
rect 1650 28696 1666 28698
rect 193 28666 219 28696
rect 1619 28666 1666 28696
rect 122 28602 188 28618
rect 122 28568 138 28602
rect 172 28600 188 28602
rect 1650 28664 1666 28666
rect 1700 28664 1716 28698
rect 1650 28648 1716 28664
rect 172 28570 219 28600
rect 1619 28570 1645 28600
rect 172 28568 188 28570
rect 122 28552 188 28568
rect 1650 28506 1716 28522
rect 1650 28504 1666 28506
rect 193 28474 219 28504
rect 1619 28474 1666 28504
rect 122 28410 188 28426
rect 122 28376 138 28410
rect 172 28408 188 28410
rect 1650 28472 1666 28474
rect 1700 28472 1716 28506
rect 1650 28456 1716 28472
rect 172 28378 219 28408
rect 1619 28378 1645 28408
rect 172 28376 188 28378
rect 122 28360 188 28376
rect 1650 28314 1716 28330
rect 1650 28312 1666 28314
rect 193 28282 219 28312
rect 1619 28282 1666 28312
rect 122 28218 188 28234
rect 122 28184 138 28218
rect 172 28216 188 28218
rect 1650 28280 1666 28282
rect 1700 28280 1716 28314
rect 1650 28264 1716 28280
rect 172 28186 219 28216
rect 1619 28186 1645 28216
rect 172 28184 188 28186
rect 122 28168 188 28184
rect 1650 28122 1716 28138
rect 1650 28120 1666 28122
rect 193 28090 219 28120
rect 1619 28090 1666 28120
rect 122 28026 188 28042
rect 122 27992 138 28026
rect 172 28024 188 28026
rect 1650 28088 1666 28090
rect 1700 28088 1716 28122
rect 1650 28072 1716 28088
rect 172 27994 219 28024
rect 1619 27994 1645 28024
rect 172 27992 188 27994
rect 122 27976 188 27992
rect 1650 27930 1716 27946
rect 1650 27928 1666 27930
rect 193 27898 219 27928
rect 1619 27898 1666 27928
rect 122 27834 188 27850
rect 122 27800 138 27834
rect 172 27832 188 27834
rect 1650 27896 1666 27898
rect 1700 27896 1716 27930
rect 1650 27880 1716 27896
rect 172 27802 219 27832
rect 1619 27802 1645 27832
rect 172 27800 188 27802
rect 122 27784 188 27800
rect 1650 27738 1716 27754
rect 1650 27736 1666 27738
rect 193 27706 219 27736
rect 1619 27706 1666 27736
rect 122 27642 188 27658
rect 122 27608 138 27642
rect 172 27640 188 27642
rect 1650 27704 1666 27706
rect 1700 27704 1716 27738
rect 1650 27688 1716 27704
rect 172 27610 219 27640
rect 1619 27610 1645 27640
rect 172 27608 188 27610
rect 122 27592 188 27608
rect 1650 27546 1716 27562
rect 1650 27544 1666 27546
rect 193 27514 219 27544
rect 1619 27514 1666 27544
rect 122 27450 188 27466
rect 122 27416 138 27450
rect 172 27448 188 27450
rect 1650 27512 1666 27514
rect 1700 27512 1716 27546
rect 1650 27496 1716 27512
rect 172 27418 219 27448
rect 1619 27418 1645 27448
rect 172 27416 188 27418
rect 122 27400 188 27416
rect 1650 27354 1716 27370
rect 1650 27352 1666 27354
rect 193 27322 219 27352
rect 1619 27322 1666 27352
rect 122 27258 188 27274
rect 122 27224 138 27258
rect 172 27256 188 27258
rect 1650 27320 1666 27322
rect 1700 27320 1716 27354
rect 1650 27304 1716 27320
rect 172 27226 219 27256
rect 1619 27226 1645 27256
rect 172 27224 188 27226
rect 122 27208 188 27224
rect 1650 27162 1716 27178
rect 1650 27160 1666 27162
rect 193 27130 219 27160
rect 1619 27130 1666 27160
rect 122 27066 188 27082
rect 122 27032 138 27066
rect 172 27064 188 27066
rect 1650 27128 1666 27130
rect 1700 27128 1716 27162
rect 1650 27112 1716 27128
rect 172 27034 219 27064
rect 1619 27034 1645 27064
rect 172 27032 188 27034
rect 122 27016 188 27032
rect 1650 26970 1716 26986
rect 1650 26968 1666 26970
rect 193 26938 219 26968
rect 1619 26938 1666 26968
rect 122 26874 188 26890
rect 122 26840 138 26874
rect 172 26872 188 26874
rect 1650 26936 1666 26938
rect 1700 26936 1716 26970
rect 1650 26920 1716 26936
rect 172 26842 219 26872
rect 1619 26842 1645 26872
rect 172 26840 188 26842
rect 122 26824 188 26840
rect 1650 26778 1716 26794
rect 1650 26776 1666 26778
rect 193 26746 219 26776
rect 1619 26746 1666 26776
rect 122 26682 188 26698
rect 122 26648 138 26682
rect 172 26680 188 26682
rect 1650 26744 1666 26746
rect 1700 26744 1716 26778
rect 1650 26728 1716 26744
rect 172 26650 219 26680
rect 1619 26650 1645 26680
rect 172 26648 188 26650
rect 122 26632 188 26648
rect 1650 26586 1716 26602
rect 1650 26584 1666 26586
rect 193 26554 219 26584
rect 1619 26554 1666 26584
rect 122 26490 188 26506
rect 122 26456 138 26490
rect 172 26488 188 26490
rect 1650 26552 1666 26554
rect 1700 26552 1716 26586
rect 1650 26536 1716 26552
rect 172 26458 219 26488
rect 1619 26458 1645 26488
rect 172 26456 188 26458
rect 122 26440 188 26456
rect 1650 26394 1716 26410
rect 1650 26392 1666 26394
rect 193 26362 219 26392
rect 1619 26362 1666 26392
rect 122 26298 188 26314
rect 122 26264 138 26298
rect 172 26296 188 26298
rect 1650 26360 1666 26362
rect 1700 26360 1716 26394
rect 1650 26344 1716 26360
rect 172 26266 219 26296
rect 1619 26266 1645 26296
rect 172 26264 188 26266
rect 122 26248 188 26264
rect 1650 26202 1716 26218
rect 1650 26200 1666 26202
rect 193 26170 219 26200
rect 1619 26170 1666 26200
rect 122 26106 188 26122
rect 122 26072 138 26106
rect 172 26104 188 26106
rect 1650 26168 1666 26170
rect 1700 26168 1716 26202
rect 1650 26152 1716 26168
rect 172 26074 219 26104
rect 1619 26074 1645 26104
rect 172 26072 188 26074
rect 122 26056 188 26072
rect 1650 26010 1716 26026
rect 1650 26008 1666 26010
rect 193 25978 219 26008
rect 1619 25978 1666 26008
rect 122 25914 188 25930
rect 122 25880 138 25914
rect 172 25912 188 25914
rect 1650 25976 1666 25978
rect 1700 25976 1716 26010
rect 1650 25960 1716 25976
rect 172 25882 219 25912
rect 1619 25882 1645 25912
rect 172 25880 188 25882
rect 122 25864 188 25880
rect 1650 25818 1716 25834
rect 1650 25816 1666 25818
rect 193 25786 219 25816
rect 1619 25786 1666 25816
rect 122 25722 188 25738
rect 122 25688 138 25722
rect 172 25720 188 25722
rect 1650 25784 1666 25786
rect 1700 25784 1716 25818
rect 1650 25768 1716 25784
rect 172 25690 219 25720
rect 1619 25690 1645 25720
rect 172 25688 188 25690
rect 122 25672 188 25688
rect 1650 25626 1716 25642
rect 1650 25624 1666 25626
rect 193 25594 219 25624
rect 1619 25594 1666 25624
rect 122 25530 188 25546
rect 122 25496 138 25530
rect 172 25528 188 25530
rect 1650 25592 1666 25594
rect 1700 25592 1716 25626
rect 1650 25576 1716 25592
rect 172 25498 219 25528
rect 1619 25498 1645 25528
rect 172 25496 188 25498
rect 122 25480 188 25496
rect 1650 25434 1716 25450
rect 1650 25432 1666 25434
rect 193 25402 219 25432
rect 1619 25402 1666 25432
rect 122 25338 188 25354
rect 122 25304 138 25338
rect 172 25336 188 25338
rect 1650 25400 1666 25402
rect 1700 25400 1716 25434
rect 1650 25384 1716 25400
rect 172 25306 219 25336
rect 1619 25306 1645 25336
rect 172 25304 188 25306
rect 122 25288 188 25304
rect 1650 25242 1716 25258
rect 1650 25240 1666 25242
rect 193 25210 219 25240
rect 1619 25210 1666 25240
rect 122 25146 188 25162
rect 122 25112 138 25146
rect 172 25144 188 25146
rect 1650 25208 1666 25210
rect 1700 25208 1716 25242
rect 1650 25192 1716 25208
rect 172 25114 219 25144
rect 1619 25114 1645 25144
rect 172 25112 188 25114
rect 122 25096 188 25112
rect 1650 25050 1716 25066
rect 1650 25048 1666 25050
rect 193 25018 219 25048
rect 1619 25018 1666 25048
rect 122 24954 188 24970
rect 122 24920 138 24954
rect 172 24952 188 24954
rect 1650 25016 1666 25018
rect 1700 25016 1716 25050
rect 1650 25000 1716 25016
rect 172 24922 219 24952
rect 1619 24922 1645 24952
rect 172 24920 188 24922
rect 122 24904 188 24920
rect 1650 24858 1716 24874
rect 1650 24856 1666 24858
rect 193 24826 219 24856
rect 1619 24826 1666 24856
rect 122 24762 188 24778
rect 122 24728 138 24762
rect 172 24760 188 24762
rect 1650 24824 1666 24826
rect 1700 24824 1716 24858
rect 1650 24808 1716 24824
rect 172 24730 219 24760
rect 1619 24730 1645 24760
rect 172 24728 188 24730
rect 122 24712 188 24728
rect 1650 24666 1716 24682
rect 1650 24664 1666 24666
rect 193 24634 219 24664
rect 1619 24634 1666 24664
rect 122 24570 188 24586
rect 122 24536 138 24570
rect 172 24568 188 24570
rect 1650 24632 1666 24634
rect 1700 24632 1716 24666
rect 1650 24616 1716 24632
rect 172 24538 219 24568
rect 1619 24538 1645 24568
rect 172 24536 188 24538
rect 122 24520 188 24536
rect 1650 24474 1716 24490
rect 1650 24472 1666 24474
rect 193 24442 219 24472
rect 1619 24442 1666 24472
rect 122 24378 188 24394
rect 122 24344 138 24378
rect 172 24376 188 24378
rect 1650 24440 1666 24442
rect 1700 24440 1716 24474
rect 1650 24424 1716 24440
rect 172 24346 219 24376
rect 1619 24346 1645 24376
rect 172 24344 188 24346
rect 122 24328 188 24344
rect 1650 24282 1716 24298
rect 1650 24280 1666 24282
rect 193 24250 219 24280
rect 1619 24250 1666 24280
rect 122 24186 188 24202
rect 122 24152 138 24186
rect 172 24184 188 24186
rect 1650 24248 1666 24250
rect 1700 24248 1716 24282
rect 1650 24232 1716 24248
rect 172 24154 219 24184
rect 1619 24154 1645 24184
rect 172 24152 188 24154
rect 122 24136 188 24152
rect 1650 24090 1716 24106
rect 1650 24088 1666 24090
rect 193 24058 219 24088
rect 1619 24058 1666 24088
rect 122 23994 188 24010
rect 122 23960 138 23994
rect 172 23992 188 23994
rect 1650 24056 1666 24058
rect 1700 24056 1716 24090
rect 1650 24040 1716 24056
rect 172 23962 219 23992
rect 1619 23962 1645 23992
rect 172 23960 188 23962
rect 122 23944 188 23960
rect 1650 23898 1716 23914
rect 1650 23896 1666 23898
rect 193 23866 219 23896
rect 1619 23866 1666 23896
rect 122 23802 188 23818
rect 122 23768 138 23802
rect 172 23800 188 23802
rect 1650 23864 1666 23866
rect 1700 23864 1716 23898
rect 1650 23848 1716 23864
rect 172 23770 219 23800
rect 1619 23770 1645 23800
rect 172 23768 188 23770
rect 122 23752 188 23768
rect 1650 23706 1716 23722
rect 1650 23704 1666 23706
rect 193 23674 219 23704
rect 1619 23674 1666 23704
rect 122 23610 188 23626
rect 122 23576 138 23610
rect 172 23608 188 23610
rect 1650 23672 1666 23674
rect 1700 23672 1716 23706
rect 1650 23656 1716 23672
rect 172 23578 219 23608
rect 1619 23578 1645 23608
rect 172 23576 188 23578
rect 122 23560 188 23576
rect 1650 23514 1716 23530
rect 1650 23512 1666 23514
rect 193 23482 219 23512
rect 1619 23482 1666 23512
rect 122 23418 188 23434
rect 122 23384 138 23418
rect 172 23416 188 23418
rect 1650 23480 1666 23482
rect 1700 23480 1716 23514
rect 1650 23464 1716 23480
rect 172 23386 219 23416
rect 1619 23386 1645 23416
rect 172 23384 188 23386
rect 122 23368 188 23384
rect 1650 23322 1716 23338
rect 1650 23320 1666 23322
rect 193 23290 219 23320
rect 1619 23290 1666 23320
rect 122 23226 188 23242
rect 122 23192 138 23226
rect 172 23224 188 23226
rect 1650 23288 1666 23290
rect 1700 23288 1716 23322
rect 1650 23272 1716 23288
rect 172 23194 219 23224
rect 1619 23194 1645 23224
rect 172 23192 188 23194
rect 122 23176 188 23192
rect 1650 23130 1716 23146
rect 1650 23128 1666 23130
rect 193 23098 219 23128
rect 1619 23098 1666 23128
rect 1650 23096 1666 23098
rect 1700 23096 1716 23130
rect 1650 23080 1716 23096
rect 122 21656 188 21672
rect 122 21622 138 21656
rect 172 21654 188 21656
rect 172 21624 219 21654
rect 1619 21624 1645 21654
rect 172 21622 188 21624
rect 122 21606 188 21622
rect 1650 21560 1716 21576
rect 1650 21558 1666 21560
rect 193 21528 219 21558
rect 1619 21528 1666 21558
rect 122 21464 188 21480
rect 122 21430 138 21464
rect 172 21462 188 21464
rect 1650 21526 1666 21528
rect 1700 21526 1716 21560
rect 1650 21510 1716 21526
rect 172 21432 219 21462
rect 1619 21432 1645 21462
rect 172 21430 188 21432
rect 122 21414 188 21430
rect 1650 21368 1716 21384
rect 1650 21366 1666 21368
rect 193 21336 219 21366
rect 1619 21336 1666 21366
rect 122 21272 188 21288
rect 122 21238 138 21272
rect 172 21270 188 21272
rect 1650 21334 1666 21336
rect 1700 21334 1716 21368
rect 1650 21318 1716 21334
rect 172 21240 219 21270
rect 1619 21240 1645 21270
rect 172 21238 188 21240
rect 122 21222 188 21238
rect 1650 21176 1716 21192
rect 1650 21174 1666 21176
rect 193 21144 219 21174
rect 1619 21144 1666 21174
rect 122 21080 188 21096
rect 122 21046 138 21080
rect 172 21078 188 21080
rect 1650 21142 1666 21144
rect 1700 21142 1716 21176
rect 1650 21126 1716 21142
rect 172 21048 219 21078
rect 1619 21048 1645 21078
rect 172 21046 188 21048
rect 122 21030 188 21046
rect 1650 20984 1716 21000
rect 1650 20982 1666 20984
rect 193 20952 219 20982
rect 1619 20952 1666 20982
rect 122 20888 188 20904
rect 122 20854 138 20888
rect 172 20886 188 20888
rect 1650 20950 1666 20952
rect 1700 20950 1716 20984
rect 1650 20934 1716 20950
rect 172 20856 219 20886
rect 1619 20856 1645 20886
rect 172 20854 188 20856
rect 122 20838 188 20854
rect 1650 20792 1716 20808
rect 1650 20790 1666 20792
rect 193 20760 219 20790
rect 1619 20760 1666 20790
rect 122 20696 188 20712
rect 122 20662 138 20696
rect 172 20694 188 20696
rect 1650 20758 1666 20760
rect 1700 20758 1716 20792
rect 1650 20742 1716 20758
rect 172 20664 219 20694
rect 1619 20664 1645 20694
rect 172 20662 188 20664
rect 122 20646 188 20662
rect 1650 20600 1716 20616
rect 1650 20598 1666 20600
rect 193 20568 219 20598
rect 1619 20568 1666 20598
rect 122 20504 188 20520
rect 122 20470 138 20504
rect 172 20502 188 20504
rect 1650 20566 1666 20568
rect 1700 20566 1716 20600
rect 1650 20550 1716 20566
rect 172 20472 219 20502
rect 1619 20472 1645 20502
rect 172 20470 188 20472
rect 122 20454 188 20470
rect 1650 20408 1716 20424
rect 1650 20406 1666 20408
rect 193 20376 219 20406
rect 1619 20376 1666 20406
rect 122 20312 188 20328
rect 122 20278 138 20312
rect 172 20310 188 20312
rect 1650 20374 1666 20376
rect 1700 20374 1716 20408
rect 1650 20358 1716 20374
rect 172 20280 219 20310
rect 1619 20280 1645 20310
rect 172 20278 188 20280
rect 122 20262 188 20278
rect 1650 20216 1716 20232
rect 1650 20214 1666 20216
rect 193 20184 219 20214
rect 1619 20184 1666 20214
rect 122 20120 188 20136
rect 122 20086 138 20120
rect 172 20118 188 20120
rect 1650 20182 1666 20184
rect 1700 20182 1716 20216
rect 1650 20166 1716 20182
rect 172 20088 219 20118
rect 1619 20088 1645 20118
rect 172 20086 188 20088
rect 122 20070 188 20086
rect 1650 20024 1716 20040
rect 1650 20022 1666 20024
rect 193 19992 219 20022
rect 1619 19992 1666 20022
rect 122 19928 188 19944
rect 122 19894 138 19928
rect 172 19926 188 19928
rect 1650 19990 1666 19992
rect 1700 19990 1716 20024
rect 1650 19974 1716 19990
rect 172 19896 219 19926
rect 1619 19896 1645 19926
rect 172 19894 188 19896
rect 122 19878 188 19894
rect 1650 19832 1716 19848
rect 1650 19830 1666 19832
rect 193 19800 219 19830
rect 1619 19800 1666 19830
rect 122 19736 188 19752
rect 122 19702 138 19736
rect 172 19734 188 19736
rect 1650 19798 1666 19800
rect 1700 19798 1716 19832
rect 1650 19782 1716 19798
rect 172 19704 219 19734
rect 1619 19704 1645 19734
rect 172 19702 188 19704
rect 122 19686 188 19702
rect 1650 19640 1716 19656
rect 1650 19638 1666 19640
rect 193 19608 219 19638
rect 1619 19608 1666 19638
rect 122 19544 188 19560
rect 122 19510 138 19544
rect 172 19542 188 19544
rect 1650 19606 1666 19608
rect 1700 19606 1716 19640
rect 1650 19590 1716 19606
rect 172 19512 219 19542
rect 1619 19512 1645 19542
rect 172 19510 188 19512
rect 122 19494 188 19510
rect 1650 19448 1716 19464
rect 1650 19446 1666 19448
rect 193 19416 219 19446
rect 1619 19416 1666 19446
rect 122 19352 188 19368
rect 122 19318 138 19352
rect 172 19350 188 19352
rect 1650 19414 1666 19416
rect 1700 19414 1716 19448
rect 1650 19398 1716 19414
rect 172 19320 219 19350
rect 1619 19320 1645 19350
rect 172 19318 188 19320
rect 122 19302 188 19318
rect 1650 19256 1716 19272
rect 1650 19254 1666 19256
rect 193 19224 219 19254
rect 1619 19224 1666 19254
rect 122 19160 188 19176
rect 122 19126 138 19160
rect 172 19158 188 19160
rect 1650 19222 1666 19224
rect 1700 19222 1716 19256
rect 1650 19206 1716 19222
rect 172 19128 219 19158
rect 1619 19128 1645 19158
rect 172 19126 188 19128
rect 122 19110 188 19126
rect 1650 19064 1716 19080
rect 1650 19062 1666 19064
rect 193 19032 219 19062
rect 1619 19032 1666 19062
rect 122 18968 188 18984
rect 122 18934 138 18968
rect 172 18966 188 18968
rect 1650 19030 1666 19032
rect 1700 19030 1716 19064
rect 1650 19014 1716 19030
rect 172 18936 219 18966
rect 1619 18936 1645 18966
rect 172 18934 188 18936
rect 122 18918 188 18934
rect 1650 18872 1716 18888
rect 1650 18870 1666 18872
rect 193 18840 219 18870
rect 1619 18840 1666 18870
rect 122 18776 188 18792
rect 122 18742 138 18776
rect 172 18774 188 18776
rect 1650 18838 1666 18840
rect 1700 18838 1716 18872
rect 1650 18822 1716 18838
rect 172 18744 219 18774
rect 1619 18744 1645 18774
rect 172 18742 188 18744
rect 122 18726 188 18742
rect 1650 18680 1716 18696
rect 1650 18678 1666 18680
rect 193 18648 219 18678
rect 1619 18648 1666 18678
rect 122 18584 188 18600
rect 122 18550 138 18584
rect 172 18582 188 18584
rect 1650 18646 1666 18648
rect 1700 18646 1716 18680
rect 1650 18630 1716 18646
rect 172 18552 219 18582
rect 1619 18552 1645 18582
rect 172 18550 188 18552
rect 122 18534 188 18550
rect 1650 18488 1716 18504
rect 1650 18486 1666 18488
rect 193 18456 219 18486
rect 1619 18456 1666 18486
rect 122 18392 188 18408
rect 122 18358 138 18392
rect 172 18390 188 18392
rect 1650 18454 1666 18456
rect 1700 18454 1716 18488
rect 1650 18438 1716 18454
rect 172 18360 219 18390
rect 1619 18360 1645 18390
rect 172 18358 188 18360
rect 122 18342 188 18358
rect 1650 18296 1716 18312
rect 1650 18294 1666 18296
rect 193 18264 219 18294
rect 1619 18264 1666 18294
rect 122 18200 188 18216
rect 122 18166 138 18200
rect 172 18198 188 18200
rect 1650 18262 1666 18264
rect 1700 18262 1716 18296
rect 1650 18246 1716 18262
rect 172 18168 219 18198
rect 1619 18168 1645 18198
rect 172 18166 188 18168
rect 122 18150 188 18166
rect 1650 18104 1716 18120
rect 1650 18102 1666 18104
rect 193 18072 219 18102
rect 1619 18072 1666 18102
rect 122 18008 188 18024
rect 122 17974 138 18008
rect 172 18006 188 18008
rect 1650 18070 1666 18072
rect 1700 18070 1716 18104
rect 1650 18054 1716 18070
rect 172 17976 219 18006
rect 1619 17976 1645 18006
rect 172 17974 188 17976
rect 122 17958 188 17974
rect 1650 17912 1716 17928
rect 1650 17910 1666 17912
rect 193 17880 219 17910
rect 1619 17880 1666 17910
rect 122 17816 188 17832
rect 122 17782 138 17816
rect 172 17814 188 17816
rect 1650 17878 1666 17880
rect 1700 17878 1716 17912
rect 1650 17862 1716 17878
rect 172 17784 219 17814
rect 1619 17784 1645 17814
rect 172 17782 188 17784
rect 122 17766 188 17782
rect 1650 17720 1716 17736
rect 1650 17718 1666 17720
rect 193 17688 219 17718
rect 1619 17688 1666 17718
rect 122 17624 188 17640
rect 122 17590 138 17624
rect 172 17622 188 17624
rect 1650 17686 1666 17688
rect 1700 17686 1716 17720
rect 1650 17670 1716 17686
rect 172 17592 219 17622
rect 1619 17592 1645 17622
rect 172 17590 188 17592
rect 122 17574 188 17590
rect 1650 17528 1716 17544
rect 1650 17526 1666 17528
rect 193 17496 219 17526
rect 1619 17496 1666 17526
rect 122 17432 188 17448
rect 122 17398 138 17432
rect 172 17430 188 17432
rect 1650 17494 1666 17496
rect 1700 17494 1716 17528
rect 1650 17478 1716 17494
rect 172 17400 219 17430
rect 1619 17400 1645 17430
rect 172 17398 188 17400
rect 122 17382 188 17398
rect 1650 17336 1716 17352
rect 1650 17334 1666 17336
rect 193 17304 219 17334
rect 1619 17304 1666 17334
rect 122 17240 188 17256
rect 122 17206 138 17240
rect 172 17238 188 17240
rect 1650 17302 1666 17304
rect 1700 17302 1716 17336
rect 1650 17286 1716 17302
rect 172 17208 219 17238
rect 1619 17208 1645 17238
rect 172 17206 188 17208
rect 122 17190 188 17206
rect 1650 17144 1716 17160
rect 1650 17142 1666 17144
rect 193 17112 219 17142
rect 1619 17112 1666 17142
rect 122 17048 188 17064
rect 122 17014 138 17048
rect 172 17046 188 17048
rect 1650 17110 1666 17112
rect 1700 17110 1716 17144
rect 1650 17094 1716 17110
rect 172 17016 219 17046
rect 1619 17016 1645 17046
rect 172 17014 188 17016
rect 122 16998 188 17014
rect 1650 16952 1716 16968
rect 1650 16950 1666 16952
rect 193 16920 219 16950
rect 1619 16920 1666 16950
rect 122 16856 188 16872
rect 122 16822 138 16856
rect 172 16854 188 16856
rect 1650 16918 1666 16920
rect 1700 16918 1716 16952
rect 1650 16902 1716 16918
rect 172 16824 219 16854
rect 1619 16824 1645 16854
rect 172 16822 188 16824
rect 122 16806 188 16822
rect 1650 16760 1716 16776
rect 1650 16758 1666 16760
rect 193 16728 219 16758
rect 1619 16728 1666 16758
rect 122 16664 188 16680
rect 122 16630 138 16664
rect 172 16662 188 16664
rect 1650 16726 1666 16728
rect 1700 16726 1716 16760
rect 1650 16710 1716 16726
rect 172 16632 219 16662
rect 1619 16632 1645 16662
rect 172 16630 188 16632
rect 122 16614 188 16630
rect 1650 16568 1716 16584
rect 1650 16566 1666 16568
rect 193 16536 219 16566
rect 1619 16536 1666 16566
rect 122 16472 188 16488
rect 122 16438 138 16472
rect 172 16470 188 16472
rect 1650 16534 1666 16536
rect 1700 16534 1716 16568
rect 1650 16518 1716 16534
rect 172 16440 219 16470
rect 1619 16440 1645 16470
rect 172 16438 188 16440
rect 122 16422 188 16438
rect 1650 16376 1716 16392
rect 1650 16374 1666 16376
rect 193 16344 219 16374
rect 1619 16344 1666 16374
rect 122 16280 188 16296
rect 122 16246 138 16280
rect 172 16278 188 16280
rect 1650 16342 1666 16344
rect 1700 16342 1716 16376
rect 1650 16326 1716 16342
rect 172 16248 219 16278
rect 1619 16248 1645 16278
rect 172 16246 188 16248
rect 122 16230 188 16246
rect 1650 16184 1716 16200
rect 1650 16182 1666 16184
rect 193 16152 219 16182
rect 1619 16152 1666 16182
rect 122 16088 188 16104
rect 122 16054 138 16088
rect 172 16086 188 16088
rect 1650 16150 1666 16152
rect 1700 16150 1716 16184
rect 1650 16134 1716 16150
rect 172 16056 219 16086
rect 1619 16056 1645 16086
rect 172 16054 188 16056
rect 122 16038 188 16054
rect 1650 15992 1716 16008
rect 1650 15990 1666 15992
rect 193 15960 219 15990
rect 1619 15960 1666 15990
rect 122 15896 188 15912
rect 122 15862 138 15896
rect 172 15894 188 15896
rect 1650 15958 1666 15960
rect 1700 15958 1716 15992
rect 1650 15942 1716 15958
rect 172 15864 219 15894
rect 1619 15864 1645 15894
rect 172 15862 188 15864
rect 122 15846 188 15862
rect 1650 15800 1716 15816
rect 1650 15798 1666 15800
rect 193 15768 219 15798
rect 1619 15768 1666 15798
rect 122 15704 188 15720
rect 122 15670 138 15704
rect 172 15702 188 15704
rect 1650 15766 1666 15768
rect 1700 15766 1716 15800
rect 1650 15750 1716 15766
rect 172 15672 219 15702
rect 1619 15672 1645 15702
rect 172 15670 188 15672
rect 122 15654 188 15670
rect 1650 15608 1716 15624
rect 1650 15606 1666 15608
rect 193 15576 219 15606
rect 1619 15576 1666 15606
rect 122 15512 188 15528
rect 122 15478 138 15512
rect 172 15510 188 15512
rect 1650 15574 1666 15576
rect 1700 15574 1716 15608
rect 1650 15558 1716 15574
rect 172 15480 219 15510
rect 1619 15480 1645 15510
rect 172 15478 188 15480
rect 122 15462 188 15478
rect 1650 15416 1716 15432
rect 1650 15414 1666 15416
rect 193 15384 219 15414
rect 1619 15384 1666 15414
rect 122 15320 188 15336
rect 122 15286 138 15320
rect 172 15318 188 15320
rect 1650 15382 1666 15384
rect 1700 15382 1716 15416
rect 1650 15366 1716 15382
rect 172 15288 219 15318
rect 1619 15288 1645 15318
rect 172 15286 188 15288
rect 122 15270 188 15286
rect 1650 15224 1716 15240
rect 1650 15222 1666 15224
rect 193 15192 219 15222
rect 1619 15192 1666 15222
rect 122 15128 188 15144
rect 122 15094 138 15128
rect 172 15126 188 15128
rect 1650 15190 1666 15192
rect 1700 15190 1716 15224
rect 1650 15174 1716 15190
rect 172 15096 219 15126
rect 1619 15096 1645 15126
rect 172 15094 188 15096
rect 122 15078 188 15094
rect 1650 15032 1716 15048
rect 1650 15030 1666 15032
rect 193 15000 219 15030
rect 1619 15000 1666 15030
rect 122 14936 188 14952
rect 122 14902 138 14936
rect 172 14934 188 14936
rect 1650 14998 1666 15000
rect 1700 14998 1716 15032
rect 1650 14982 1716 14998
rect 172 14904 219 14934
rect 1619 14904 1645 14934
rect 172 14902 188 14904
rect 122 14886 188 14902
rect 1650 14840 1716 14856
rect 1650 14838 1666 14840
rect 193 14808 219 14838
rect 1619 14808 1666 14838
rect 122 14744 188 14760
rect 122 14710 138 14744
rect 172 14742 188 14744
rect 1650 14806 1666 14808
rect 1700 14806 1716 14840
rect 1650 14790 1716 14806
rect 172 14712 219 14742
rect 1619 14712 1645 14742
rect 172 14710 188 14712
rect 122 14694 188 14710
rect 1650 14648 1716 14664
rect 1650 14646 1666 14648
rect 193 14616 219 14646
rect 1619 14616 1666 14646
rect 122 14552 188 14568
rect 122 14518 138 14552
rect 172 14550 188 14552
rect 1650 14614 1666 14616
rect 1700 14614 1716 14648
rect 1650 14598 1716 14614
rect 172 14520 219 14550
rect 1619 14520 1645 14550
rect 172 14518 188 14520
rect 122 14502 188 14518
rect 1650 14456 1716 14472
rect 1650 14454 1666 14456
rect 193 14424 219 14454
rect 1619 14424 1666 14454
rect 122 14360 188 14376
rect 122 14326 138 14360
rect 172 14358 188 14360
rect 1650 14422 1666 14424
rect 1700 14422 1716 14456
rect 1650 14406 1716 14422
rect 172 14328 219 14358
rect 1619 14328 1645 14358
rect 172 14326 188 14328
rect 122 14310 188 14326
rect 1650 14264 1716 14280
rect 1650 14262 1666 14264
rect 193 14232 219 14262
rect 1619 14232 1666 14262
rect 122 14168 188 14184
rect 122 14134 138 14168
rect 172 14166 188 14168
rect 1650 14230 1666 14232
rect 1700 14230 1716 14264
rect 1650 14214 1716 14230
rect 172 14136 219 14166
rect 1619 14136 1645 14166
rect 172 14134 188 14136
rect 122 14118 188 14134
rect 1650 14072 1716 14088
rect 1650 14070 1666 14072
rect 193 14040 219 14070
rect 1619 14040 1666 14070
rect 122 13976 188 13992
rect 122 13942 138 13976
rect 172 13974 188 13976
rect 1650 14038 1666 14040
rect 1700 14038 1716 14072
rect 1650 14022 1716 14038
rect 172 13944 219 13974
rect 1619 13944 1645 13974
rect 172 13942 188 13944
rect 122 13926 188 13942
rect 1650 13880 1716 13896
rect 1650 13878 1666 13880
rect 193 13848 219 13878
rect 1619 13848 1666 13878
rect 122 13784 188 13800
rect 122 13750 138 13784
rect 172 13782 188 13784
rect 1650 13846 1666 13848
rect 1700 13846 1716 13880
rect 1650 13830 1716 13846
rect 172 13752 219 13782
rect 1619 13752 1645 13782
rect 172 13750 188 13752
rect 122 13734 188 13750
rect 1650 13688 1716 13704
rect 1650 13686 1666 13688
rect 193 13656 219 13686
rect 1619 13656 1666 13686
rect 122 13592 188 13608
rect 122 13558 138 13592
rect 172 13590 188 13592
rect 1650 13654 1666 13656
rect 1700 13654 1716 13688
rect 1650 13638 1716 13654
rect 172 13560 219 13590
rect 1619 13560 1645 13590
rect 172 13558 188 13560
rect 122 13542 188 13558
rect 1650 13496 1716 13512
rect 1650 13494 1666 13496
rect 193 13464 219 13494
rect 1619 13464 1666 13494
rect 122 13400 188 13416
rect 122 13366 138 13400
rect 172 13398 188 13400
rect 1650 13462 1666 13464
rect 1700 13462 1716 13496
rect 1650 13446 1716 13462
rect 172 13368 219 13398
rect 1619 13368 1645 13398
rect 172 13366 188 13368
rect 122 13350 188 13366
rect 1650 13304 1716 13320
rect 1650 13302 1666 13304
rect 193 13272 219 13302
rect 1619 13272 1666 13302
rect 122 13208 188 13224
rect 122 13174 138 13208
rect 172 13206 188 13208
rect 1650 13270 1666 13272
rect 1700 13270 1716 13304
rect 1650 13254 1716 13270
rect 172 13176 219 13206
rect 1619 13176 1645 13206
rect 172 13174 188 13176
rect 122 13158 188 13174
rect 1650 13112 1716 13128
rect 1650 13110 1666 13112
rect 193 13080 219 13110
rect 1619 13080 1666 13110
rect 122 13016 188 13032
rect 122 12982 138 13016
rect 172 13014 188 13016
rect 1650 13078 1666 13080
rect 1700 13078 1716 13112
rect 1650 13062 1716 13078
rect 172 12984 219 13014
rect 1619 12984 1645 13014
rect 172 12982 188 12984
rect 122 12966 188 12982
rect 1650 12920 1716 12936
rect 1650 12918 1666 12920
rect 193 12888 219 12918
rect 1619 12888 1666 12918
rect 122 12824 188 12840
rect 122 12790 138 12824
rect 172 12822 188 12824
rect 1650 12886 1666 12888
rect 1700 12886 1716 12920
rect 1650 12870 1716 12886
rect 172 12792 219 12822
rect 1619 12792 1645 12822
rect 172 12790 188 12792
rect 122 12774 188 12790
rect 1650 12728 1716 12744
rect 1650 12726 1666 12728
rect 193 12696 219 12726
rect 1619 12696 1666 12726
rect 122 12632 188 12648
rect 122 12598 138 12632
rect 172 12630 188 12632
rect 1650 12694 1666 12696
rect 1700 12694 1716 12728
rect 1650 12678 1716 12694
rect 172 12600 219 12630
rect 1619 12600 1645 12630
rect 172 12598 188 12600
rect 122 12582 188 12598
rect 1650 12536 1716 12552
rect 1650 12534 1666 12536
rect 193 12504 219 12534
rect 1619 12504 1666 12534
rect 122 12440 188 12456
rect 122 12406 138 12440
rect 172 12438 188 12440
rect 1650 12502 1666 12504
rect 1700 12502 1716 12536
rect 1650 12486 1716 12502
rect 172 12408 219 12438
rect 1619 12408 1645 12438
rect 172 12406 188 12408
rect 122 12390 188 12406
rect 1650 12344 1716 12360
rect 1650 12342 1666 12344
rect 193 12312 219 12342
rect 1619 12312 1666 12342
rect 122 12248 188 12264
rect 122 12214 138 12248
rect 172 12246 188 12248
rect 1650 12310 1666 12312
rect 1700 12310 1716 12344
rect 1650 12294 1716 12310
rect 172 12216 219 12246
rect 1619 12216 1645 12246
rect 172 12214 188 12216
rect 122 12198 188 12214
rect 1650 12152 1716 12168
rect 1650 12150 1666 12152
rect 193 12120 219 12150
rect 1619 12120 1666 12150
rect 122 12056 188 12072
rect 122 12022 138 12056
rect 172 12054 188 12056
rect 1650 12118 1666 12120
rect 1700 12118 1716 12152
rect 1650 12102 1716 12118
rect 172 12024 219 12054
rect 1619 12024 1645 12054
rect 172 12022 188 12024
rect 122 12006 188 12022
rect 1650 11960 1716 11976
rect 1650 11958 1666 11960
rect 193 11928 219 11958
rect 1619 11928 1666 11958
rect 122 11864 188 11880
rect 122 11830 138 11864
rect 172 11862 188 11864
rect 1650 11926 1666 11928
rect 1700 11926 1716 11960
rect 1650 11910 1716 11926
rect 172 11832 219 11862
rect 1619 11832 1645 11862
rect 172 11830 188 11832
rect 122 11814 188 11830
rect 1650 11768 1716 11784
rect 1650 11766 1666 11768
rect 193 11736 219 11766
rect 1619 11736 1666 11766
rect 122 11672 188 11688
rect 122 11638 138 11672
rect 172 11670 188 11672
rect 1650 11734 1666 11736
rect 1700 11734 1716 11768
rect 1650 11718 1716 11734
rect 172 11640 219 11670
rect 1619 11640 1645 11670
rect 172 11638 188 11640
rect 122 11622 188 11638
rect 1650 11576 1716 11592
rect 1650 11574 1666 11576
rect 193 11544 219 11574
rect 1619 11544 1666 11574
rect 122 11480 188 11496
rect 122 11446 138 11480
rect 172 11478 188 11480
rect 1650 11542 1666 11544
rect 1700 11542 1716 11576
rect 1650 11526 1716 11542
rect 172 11448 219 11478
rect 1619 11448 1645 11478
rect 172 11446 188 11448
rect 122 11430 188 11446
rect 1650 11384 1716 11400
rect 1650 11382 1666 11384
rect 193 11352 219 11382
rect 1619 11352 1666 11382
rect 122 11288 188 11304
rect 122 11254 138 11288
rect 172 11286 188 11288
rect 1650 11350 1666 11352
rect 1700 11350 1716 11384
rect 1650 11334 1716 11350
rect 172 11256 219 11286
rect 1619 11256 1645 11286
rect 172 11254 188 11256
rect 122 11238 188 11254
rect 1650 11192 1716 11208
rect 1650 11190 1666 11192
rect 193 11160 219 11190
rect 1619 11160 1666 11190
rect 122 11096 188 11112
rect 122 11062 138 11096
rect 172 11094 188 11096
rect 1650 11158 1666 11160
rect 1700 11158 1716 11192
rect 1650 11142 1716 11158
rect 172 11064 219 11094
rect 1619 11064 1645 11094
rect 172 11062 188 11064
rect 122 11046 188 11062
rect 1650 11000 1716 11016
rect 1650 10998 1666 11000
rect 193 10968 219 10998
rect 1619 10968 1666 10998
rect 122 10904 188 10920
rect 122 10870 138 10904
rect 172 10902 188 10904
rect 1650 10966 1666 10968
rect 1700 10966 1716 11000
rect 1650 10950 1716 10966
rect 172 10872 219 10902
rect 1619 10872 1645 10902
rect 172 10870 188 10872
rect 122 10854 188 10870
rect 1650 10808 1716 10824
rect 1650 10806 1666 10808
rect 193 10776 219 10806
rect 1619 10776 1666 10806
rect 122 10712 188 10728
rect 122 10678 138 10712
rect 172 10710 188 10712
rect 1650 10774 1666 10776
rect 1700 10774 1716 10808
rect 1650 10758 1716 10774
rect 172 10680 219 10710
rect 1619 10680 1645 10710
rect 172 10678 188 10680
rect 122 10662 188 10678
rect 1650 10616 1716 10632
rect 1650 10614 1666 10616
rect 193 10584 219 10614
rect 1619 10584 1666 10614
rect 122 10520 188 10536
rect 122 10486 138 10520
rect 172 10518 188 10520
rect 1650 10582 1666 10584
rect 1700 10582 1716 10616
rect 1650 10566 1716 10582
rect 172 10488 219 10518
rect 1619 10488 1645 10518
rect 172 10486 188 10488
rect 122 10470 188 10486
rect 1650 10424 1716 10440
rect 1650 10422 1666 10424
rect 193 10392 219 10422
rect 1619 10392 1666 10422
rect 122 10328 188 10344
rect 122 10294 138 10328
rect 172 10326 188 10328
rect 1650 10390 1666 10392
rect 1700 10390 1716 10424
rect 1650 10374 1716 10390
rect 172 10296 219 10326
rect 1619 10296 1645 10326
rect 172 10294 188 10296
rect 122 10278 188 10294
rect 1650 10232 1716 10248
rect 1650 10230 1666 10232
rect 193 10200 219 10230
rect 1619 10200 1666 10230
rect 122 10136 188 10152
rect 122 10102 138 10136
rect 172 10134 188 10136
rect 1650 10198 1666 10200
rect 1700 10198 1716 10232
rect 1650 10182 1716 10198
rect 172 10104 219 10134
rect 1619 10104 1645 10134
rect 172 10102 188 10104
rect 122 10086 188 10102
rect 1650 10040 1716 10056
rect 1650 10038 1666 10040
rect 193 10008 219 10038
rect 1619 10008 1666 10038
rect 122 9944 188 9960
rect 122 9910 138 9944
rect 172 9942 188 9944
rect 1650 10006 1666 10008
rect 1700 10006 1716 10040
rect 1650 9990 1716 10006
rect 172 9912 219 9942
rect 1619 9912 1645 9942
rect 172 9910 188 9912
rect 122 9894 188 9910
rect 1650 9848 1716 9864
rect 1650 9846 1666 9848
rect 193 9816 219 9846
rect 1619 9816 1666 9846
rect 122 9752 188 9768
rect 122 9718 138 9752
rect 172 9750 188 9752
rect 1650 9814 1666 9816
rect 1700 9814 1716 9848
rect 1650 9798 1716 9814
rect 172 9720 219 9750
rect 1619 9720 1645 9750
rect 172 9718 188 9720
rect 122 9702 188 9718
rect 1650 9656 1716 9672
rect 1650 9654 1666 9656
rect 193 9624 219 9654
rect 1619 9624 1666 9654
rect 122 9560 188 9576
rect 122 9526 138 9560
rect 172 9558 188 9560
rect 1650 9622 1666 9624
rect 1700 9622 1716 9656
rect 1650 9606 1716 9622
rect 172 9528 219 9558
rect 1619 9528 1645 9558
rect 172 9526 188 9528
rect 122 9510 188 9526
rect 1650 9464 1716 9480
rect 1650 9462 1666 9464
rect 193 9432 219 9462
rect 1619 9432 1666 9462
rect 122 9368 188 9384
rect 122 9334 138 9368
rect 172 9366 188 9368
rect 1650 9430 1666 9432
rect 1700 9430 1716 9464
rect 1650 9414 1716 9430
rect 172 9336 219 9366
rect 1619 9336 1645 9366
rect 172 9334 188 9336
rect 122 9318 188 9334
rect 1650 9272 1716 9288
rect 1650 9270 1666 9272
rect 193 9240 219 9270
rect 1619 9240 1666 9270
rect 122 9176 188 9192
rect 122 9142 138 9176
rect 172 9174 188 9176
rect 1650 9238 1666 9240
rect 1700 9238 1716 9272
rect 1650 9222 1716 9238
rect 172 9144 219 9174
rect 1619 9144 1645 9174
rect 172 9142 188 9144
rect 122 9126 188 9142
rect 1650 9080 1716 9096
rect 1650 9078 1666 9080
rect 193 9048 219 9078
rect 1619 9048 1666 9078
rect 122 8984 188 9000
rect 122 8950 138 8984
rect 172 8982 188 8984
rect 1650 9046 1666 9048
rect 1700 9046 1716 9080
rect 1650 9030 1716 9046
rect 172 8952 219 8982
rect 1619 8952 1645 8982
rect 172 8950 188 8952
rect 122 8934 188 8950
rect 1650 8888 1716 8904
rect 1650 8886 1666 8888
rect 193 8856 219 8886
rect 1619 8856 1666 8886
rect 122 8792 188 8808
rect 122 8758 138 8792
rect 172 8790 188 8792
rect 1650 8854 1666 8856
rect 1700 8854 1716 8888
rect 1650 8838 1716 8854
rect 172 8760 219 8790
rect 1619 8760 1645 8790
rect 172 8758 188 8760
rect 122 8742 188 8758
rect 1650 8696 1716 8712
rect 1650 8694 1666 8696
rect 193 8664 219 8694
rect 1619 8664 1666 8694
rect 122 8600 188 8616
rect 122 8566 138 8600
rect 172 8598 188 8600
rect 1650 8662 1666 8664
rect 1700 8662 1716 8696
rect 1650 8646 1716 8662
rect 172 8568 219 8598
rect 1619 8568 1645 8598
rect 172 8566 188 8568
rect 122 8550 188 8566
rect 1650 8504 1716 8520
rect 1650 8502 1666 8504
rect 193 8472 219 8502
rect 1619 8472 1666 8502
rect 122 8408 188 8424
rect 122 8374 138 8408
rect 172 8406 188 8408
rect 1650 8470 1666 8472
rect 1700 8470 1716 8504
rect 1650 8454 1716 8470
rect 172 8376 219 8406
rect 1619 8376 1645 8406
rect 172 8374 188 8376
rect 122 8358 188 8374
rect 1650 8312 1716 8328
rect 1650 8310 1666 8312
rect 193 8280 219 8310
rect 1619 8280 1666 8310
rect 122 8216 188 8232
rect 122 8182 138 8216
rect 172 8214 188 8216
rect 1650 8278 1666 8280
rect 1700 8278 1716 8312
rect 1650 8262 1716 8278
rect 172 8184 219 8214
rect 1619 8184 1645 8214
rect 172 8182 188 8184
rect 122 8166 188 8182
rect 1650 8120 1716 8136
rect 1650 8118 1666 8120
rect 193 8088 219 8118
rect 1619 8088 1666 8118
rect 122 8024 188 8040
rect 122 7990 138 8024
rect 172 8022 188 8024
rect 1650 8086 1666 8088
rect 1700 8086 1716 8120
rect 1650 8070 1716 8086
rect 172 7992 219 8022
rect 1619 7992 1645 8022
rect 172 7990 188 7992
rect 122 7974 188 7990
rect 1650 7928 1716 7944
rect 1650 7926 1666 7928
rect 193 7896 219 7926
rect 1619 7896 1666 7926
rect 122 7832 188 7848
rect 122 7798 138 7832
rect 172 7830 188 7832
rect 1650 7894 1666 7896
rect 1700 7894 1716 7928
rect 1650 7878 1716 7894
rect 172 7800 219 7830
rect 1619 7800 1645 7830
rect 172 7798 188 7800
rect 122 7782 188 7798
rect 1650 7736 1716 7752
rect 1650 7734 1666 7736
rect 193 7704 219 7734
rect 1619 7704 1666 7734
rect 122 7640 188 7656
rect 122 7606 138 7640
rect 172 7638 188 7640
rect 1650 7702 1666 7704
rect 1700 7702 1716 7736
rect 1650 7686 1716 7702
rect 172 7608 219 7638
rect 1619 7608 1645 7638
rect 172 7606 188 7608
rect 122 7590 188 7606
rect 1650 7544 1716 7560
rect 1650 7542 1666 7544
rect 193 7512 219 7542
rect 1619 7512 1666 7542
rect 122 7448 188 7464
rect 122 7414 138 7448
rect 172 7446 188 7448
rect 1650 7510 1666 7512
rect 1700 7510 1716 7544
rect 1650 7494 1716 7510
rect 172 7416 219 7446
rect 1619 7416 1645 7446
rect 172 7414 188 7416
rect 122 7398 188 7414
rect 1650 7352 1716 7368
rect 1650 7350 1666 7352
rect 193 7320 219 7350
rect 1619 7320 1666 7350
rect 122 7256 188 7272
rect 122 7222 138 7256
rect 172 7254 188 7256
rect 1650 7318 1666 7320
rect 1700 7318 1716 7352
rect 1650 7302 1716 7318
rect 172 7224 219 7254
rect 1619 7224 1645 7254
rect 172 7222 188 7224
rect 122 7206 188 7222
rect 1650 7160 1716 7176
rect 1650 7158 1666 7160
rect 193 7128 219 7158
rect 1619 7128 1666 7158
rect 122 7064 188 7080
rect 122 7030 138 7064
rect 172 7062 188 7064
rect 1650 7126 1666 7128
rect 1700 7126 1716 7160
rect 1650 7110 1716 7126
rect 172 7032 219 7062
rect 1619 7032 1645 7062
rect 172 7030 188 7032
rect 122 7014 188 7030
rect 1650 6968 1716 6984
rect 1650 6966 1666 6968
rect 193 6936 219 6966
rect 1619 6936 1666 6966
rect 122 6872 188 6888
rect 122 6838 138 6872
rect 172 6870 188 6872
rect 1650 6934 1666 6936
rect 1700 6934 1716 6968
rect 1650 6918 1716 6934
rect 172 6840 219 6870
rect 1619 6840 1645 6870
rect 172 6838 188 6840
rect 122 6822 188 6838
rect 1650 6776 1716 6792
rect 1650 6774 1666 6776
rect 193 6744 219 6774
rect 1619 6744 1666 6774
rect 122 6680 188 6696
rect 122 6646 138 6680
rect 172 6678 188 6680
rect 1650 6742 1666 6744
rect 1700 6742 1716 6776
rect 1650 6726 1716 6742
rect 172 6648 219 6678
rect 1619 6648 1645 6678
rect 172 6646 188 6648
rect 122 6630 188 6646
rect 1650 6584 1716 6600
rect 1650 6582 1666 6584
rect 193 6552 219 6582
rect 1619 6552 1666 6582
rect 122 6488 188 6504
rect 122 6454 138 6488
rect 172 6486 188 6488
rect 1650 6550 1666 6552
rect 1700 6550 1716 6584
rect 1650 6534 1716 6550
rect 172 6456 219 6486
rect 1619 6456 1645 6486
rect 172 6454 188 6456
rect 122 6438 188 6454
rect 1650 6392 1716 6408
rect 1650 6390 1666 6392
rect 193 6360 219 6390
rect 1619 6360 1666 6390
rect 122 6296 188 6312
rect 122 6262 138 6296
rect 172 6294 188 6296
rect 1650 6358 1666 6360
rect 1700 6358 1716 6392
rect 1650 6342 1716 6358
rect 172 6264 219 6294
rect 1619 6264 1645 6294
rect 172 6262 188 6264
rect 122 6246 188 6262
rect 1650 6200 1716 6216
rect 1650 6198 1666 6200
rect 193 6168 219 6198
rect 1619 6168 1666 6198
rect 122 6104 188 6120
rect 122 6070 138 6104
rect 172 6102 188 6104
rect 1650 6166 1666 6168
rect 1700 6166 1716 6200
rect 1650 6150 1716 6166
rect 172 6072 219 6102
rect 1619 6072 1645 6102
rect 172 6070 188 6072
rect 122 6054 188 6070
rect 1650 6008 1716 6024
rect 1650 6006 1666 6008
rect 193 5976 219 6006
rect 1619 5976 1666 6006
rect 122 5912 188 5928
rect 122 5878 138 5912
rect 172 5910 188 5912
rect 1650 5974 1666 5976
rect 1700 5974 1716 6008
rect 1650 5958 1716 5974
rect 172 5880 219 5910
rect 1619 5880 1645 5910
rect 172 5878 188 5880
rect 122 5862 188 5878
rect 1650 5816 1716 5832
rect 1650 5814 1666 5816
rect 193 5784 219 5814
rect 1619 5784 1666 5814
rect 122 5720 188 5736
rect 122 5686 138 5720
rect 172 5718 188 5720
rect 1650 5782 1666 5784
rect 1700 5782 1716 5816
rect 1650 5766 1716 5782
rect 172 5688 219 5718
rect 1619 5688 1645 5718
rect 172 5686 188 5688
rect 122 5670 188 5686
rect 1650 5624 1716 5640
rect 1650 5622 1666 5624
rect 193 5592 219 5622
rect 1619 5592 1666 5622
rect 122 5528 188 5544
rect 122 5494 138 5528
rect 172 5526 188 5528
rect 1650 5590 1666 5592
rect 1700 5590 1716 5624
rect 1650 5574 1716 5590
rect 172 5496 219 5526
rect 1619 5496 1645 5526
rect 172 5494 188 5496
rect 122 5478 188 5494
rect 1650 5432 1716 5448
rect 1650 5430 1666 5432
rect 193 5400 219 5430
rect 1619 5400 1666 5430
rect 122 5336 188 5352
rect 122 5302 138 5336
rect 172 5334 188 5336
rect 1650 5398 1666 5400
rect 1700 5398 1716 5432
rect 1650 5382 1716 5398
rect 172 5304 219 5334
rect 1619 5304 1645 5334
rect 172 5302 188 5304
rect 122 5286 188 5302
rect 1650 5240 1716 5256
rect 1650 5238 1666 5240
rect 193 5208 219 5238
rect 1619 5208 1666 5238
rect 122 5144 188 5160
rect 122 5110 138 5144
rect 172 5142 188 5144
rect 1650 5206 1666 5208
rect 1700 5206 1716 5240
rect 1650 5190 1716 5206
rect 172 5112 219 5142
rect 1619 5112 1645 5142
rect 172 5110 188 5112
rect 122 5094 188 5110
rect 1650 5048 1716 5064
rect 1650 5046 1666 5048
rect 193 5016 219 5046
rect 1619 5016 1666 5046
rect 122 4952 188 4968
rect 122 4918 138 4952
rect 172 4950 188 4952
rect 1650 5014 1666 5016
rect 1700 5014 1716 5048
rect 1650 4998 1716 5014
rect 172 4920 219 4950
rect 1619 4920 1645 4950
rect 172 4918 188 4920
rect 122 4902 188 4918
rect 1650 4856 1716 4872
rect 1650 4854 1666 4856
rect 193 4824 219 4854
rect 1619 4824 1666 4854
rect 122 4760 188 4776
rect 122 4726 138 4760
rect 172 4758 188 4760
rect 1650 4822 1666 4824
rect 1700 4822 1716 4856
rect 1650 4806 1716 4822
rect 172 4728 219 4758
rect 1619 4728 1645 4758
rect 172 4726 188 4728
rect 122 4710 188 4726
rect 1650 4664 1716 4680
rect 1650 4662 1666 4664
rect 193 4632 219 4662
rect 1619 4632 1666 4662
rect 122 4568 188 4584
rect 122 4534 138 4568
rect 172 4566 188 4568
rect 1650 4630 1666 4632
rect 1700 4630 1716 4664
rect 1650 4614 1716 4630
rect 172 4536 219 4566
rect 1619 4536 1645 4566
rect 172 4534 188 4536
rect 122 4518 188 4534
rect 1650 4472 1716 4488
rect 1650 4470 1666 4472
rect 193 4440 219 4470
rect 1619 4440 1666 4470
rect 122 4376 188 4392
rect 122 4342 138 4376
rect 172 4374 188 4376
rect 1650 4438 1666 4440
rect 1700 4438 1716 4472
rect 1650 4422 1716 4438
rect 172 4344 219 4374
rect 1619 4344 1645 4374
rect 172 4342 188 4344
rect 122 4326 188 4342
rect 1650 4280 1716 4296
rect 1650 4278 1666 4280
rect 193 4248 219 4278
rect 1619 4248 1666 4278
rect 122 4184 188 4200
rect 122 4150 138 4184
rect 172 4182 188 4184
rect 1650 4246 1666 4248
rect 1700 4246 1716 4280
rect 1650 4230 1716 4246
rect 172 4152 219 4182
rect 1619 4152 1645 4182
rect 172 4150 188 4152
rect 122 4134 188 4150
rect 1650 4088 1716 4104
rect 1650 4086 1666 4088
rect 193 4056 219 4086
rect 1619 4056 1666 4086
rect 122 3992 188 4008
rect 122 3958 138 3992
rect 172 3990 188 3992
rect 1650 4054 1666 4056
rect 1700 4054 1716 4088
rect 1650 4038 1716 4054
rect 172 3960 219 3990
rect 1619 3960 1645 3990
rect 172 3958 188 3960
rect 122 3942 188 3958
rect 1650 3896 1716 3912
rect 1650 3894 1666 3896
rect 193 3864 219 3894
rect 1619 3864 1666 3894
rect 122 3800 188 3816
rect 122 3766 138 3800
rect 172 3798 188 3800
rect 1650 3862 1666 3864
rect 1700 3862 1716 3896
rect 1650 3846 1716 3862
rect 172 3768 219 3798
rect 1619 3768 1645 3798
rect 172 3766 188 3768
rect 122 3750 188 3766
rect 1650 3704 1716 3720
rect 1650 3702 1666 3704
rect 193 3672 219 3702
rect 1619 3672 1666 3702
rect 122 3608 188 3624
rect 122 3574 138 3608
rect 172 3606 188 3608
rect 1650 3670 1666 3672
rect 1700 3670 1716 3704
rect 1650 3654 1716 3670
rect 172 3576 219 3606
rect 1619 3576 1645 3606
rect 172 3574 188 3576
rect 122 3558 188 3574
rect 1650 3512 1716 3528
rect 1650 3510 1666 3512
rect 193 3480 219 3510
rect 1619 3480 1666 3510
rect 122 3416 188 3432
rect 122 3382 138 3416
rect 172 3414 188 3416
rect 1650 3478 1666 3480
rect 1700 3478 1716 3512
rect 1650 3462 1716 3478
rect 172 3384 219 3414
rect 1619 3384 1645 3414
rect 172 3382 188 3384
rect 122 3366 188 3382
rect 1650 3320 1716 3336
rect 1650 3318 1666 3320
rect 193 3288 219 3318
rect 1619 3288 1666 3318
rect 122 3224 188 3240
rect 122 3190 138 3224
rect 172 3222 188 3224
rect 1650 3286 1666 3288
rect 1700 3286 1716 3320
rect 1650 3270 1716 3286
rect 172 3192 219 3222
rect 1619 3192 1645 3222
rect 172 3190 188 3192
rect 122 3174 188 3190
rect 1650 3128 1716 3144
rect 1650 3126 1666 3128
rect 193 3096 219 3126
rect 1619 3096 1666 3126
rect 122 3032 188 3048
rect 122 2998 138 3032
rect 172 3030 188 3032
rect 1650 3094 1666 3096
rect 1700 3094 1716 3128
rect 1650 3078 1716 3094
rect 172 3000 219 3030
rect 1619 3000 1645 3030
rect 172 2998 188 3000
rect 122 2982 188 2998
rect 1650 2936 1716 2952
rect 1650 2934 1666 2936
rect 193 2904 219 2934
rect 1619 2904 1666 2934
rect 122 2840 188 2856
rect 122 2806 138 2840
rect 172 2838 188 2840
rect 1650 2902 1666 2904
rect 1700 2902 1716 2936
rect 1650 2886 1716 2902
rect 172 2808 219 2838
rect 1619 2808 1645 2838
rect 172 2806 188 2808
rect 122 2790 188 2806
rect 1650 2744 1716 2760
rect 1650 2742 1666 2744
rect 193 2712 219 2742
rect 1619 2712 1666 2742
rect 122 2648 188 2664
rect 122 2614 138 2648
rect 172 2646 188 2648
rect 1650 2710 1666 2712
rect 1700 2710 1716 2744
rect 1650 2694 1716 2710
rect 172 2616 219 2646
rect 1619 2616 1645 2646
rect 172 2614 188 2616
rect 122 2598 188 2614
rect 1650 2552 1716 2568
rect 1650 2550 1666 2552
rect 193 2520 219 2550
rect 1619 2520 1666 2550
rect 122 2456 188 2472
rect 122 2422 138 2456
rect 172 2454 188 2456
rect 1650 2518 1666 2520
rect 1700 2518 1716 2552
rect 1650 2502 1716 2518
rect 172 2424 219 2454
rect 1619 2424 1645 2454
rect 172 2422 188 2424
rect 122 2406 188 2422
rect 1650 2360 1716 2376
rect 1650 2358 1666 2360
rect 193 2328 219 2358
rect 1619 2328 1666 2358
rect 122 2264 188 2280
rect 122 2230 138 2264
rect 172 2262 188 2264
rect 1650 2326 1666 2328
rect 1700 2326 1716 2360
rect 1650 2310 1716 2326
rect 172 2232 219 2262
rect 1619 2232 1645 2262
rect 172 2230 188 2232
rect 122 2214 188 2230
rect 1650 2168 1716 2184
rect 1650 2166 1666 2168
rect 193 2136 219 2166
rect 1619 2136 1666 2166
rect 122 2072 188 2088
rect 122 2038 138 2072
rect 172 2070 188 2072
rect 1650 2134 1666 2136
rect 1700 2134 1716 2168
rect 1650 2118 1716 2134
rect 172 2040 219 2070
rect 1619 2040 1645 2070
rect 172 2038 188 2040
rect 122 2022 188 2038
rect 1650 1976 1716 1992
rect 1650 1974 1666 1976
rect 193 1944 219 1974
rect 1619 1944 1666 1974
rect 122 1880 188 1896
rect 122 1846 138 1880
rect 172 1878 188 1880
rect 1650 1942 1666 1944
rect 1700 1942 1716 1976
rect 1650 1926 1716 1942
rect 172 1848 219 1878
rect 1619 1848 1645 1878
rect 172 1846 188 1848
rect 122 1830 188 1846
rect 1650 1784 1716 1800
rect 1650 1782 1666 1784
rect 193 1752 219 1782
rect 1619 1752 1666 1782
rect 122 1688 188 1704
rect 122 1654 138 1688
rect 172 1686 188 1688
rect 1650 1750 1666 1752
rect 1700 1750 1716 1784
rect 1650 1734 1716 1750
rect 172 1656 219 1686
rect 1619 1656 1645 1686
rect 172 1654 188 1656
rect 122 1638 188 1654
rect 1650 1592 1716 1608
rect 1650 1590 1666 1592
rect 193 1560 219 1590
rect 1619 1560 1666 1590
rect 122 1496 188 1512
rect 122 1462 138 1496
rect 172 1494 188 1496
rect 1650 1558 1666 1560
rect 1700 1558 1716 1592
rect 1650 1542 1716 1558
rect 172 1464 219 1494
rect 1619 1464 1645 1494
rect 172 1462 188 1464
rect 122 1446 188 1462
rect 1650 1400 1716 1416
rect 1650 1398 1666 1400
rect 193 1368 219 1398
rect 1619 1368 1666 1398
rect 122 1304 188 1320
rect 122 1270 138 1304
rect 172 1302 188 1304
rect 1650 1366 1666 1368
rect 1700 1366 1716 1400
rect 1650 1350 1716 1366
rect 172 1272 219 1302
rect 1619 1272 1645 1302
rect 172 1270 188 1272
rect 122 1254 188 1270
rect 1650 1208 1716 1224
rect 1650 1206 1666 1208
rect 193 1176 219 1206
rect 1619 1176 1666 1206
rect 122 1112 188 1128
rect 122 1078 138 1112
rect 172 1110 188 1112
rect 1650 1174 1666 1176
rect 1700 1174 1716 1208
rect 1650 1158 1716 1174
rect 172 1080 219 1110
rect 1619 1080 1645 1110
rect 172 1078 188 1080
rect 122 1062 188 1078
rect 1650 1016 1716 1032
rect 1650 1014 1666 1016
rect 193 984 219 1014
rect 1619 984 1666 1014
rect 122 920 188 936
rect 122 886 138 920
rect 172 918 188 920
rect 1650 982 1666 984
rect 1700 982 1716 1016
rect 1650 966 1716 982
rect 172 888 219 918
rect 1619 888 1645 918
rect 172 886 188 888
rect 122 870 188 886
rect 1650 824 1716 840
rect 1650 822 1666 824
rect 193 792 219 822
rect 1619 792 1666 822
rect 122 728 188 744
rect 122 694 138 728
rect 172 726 188 728
rect 1650 790 1666 792
rect 1700 790 1716 824
rect 1650 774 1716 790
rect 172 696 219 726
rect 1619 696 1645 726
rect 172 694 188 696
rect 122 678 188 694
rect 1650 632 1716 648
rect 1650 630 1666 632
rect 193 600 219 630
rect 1619 600 1666 630
rect 1650 598 1666 600
rect 1700 598 1716 632
rect 1650 582 1716 598
<< polycont >>
rect 138 44120 172 44154
rect 138 43928 172 43962
rect 1666 44024 1700 44058
rect 138 43736 172 43770
rect 1666 43832 1700 43866
rect 138 43544 172 43578
rect 1666 43640 1700 43674
rect 138 43352 172 43386
rect 1666 43448 1700 43482
rect 138 43160 172 43194
rect 1666 43256 1700 43290
rect 138 42968 172 43002
rect 1666 43064 1700 43098
rect 138 42776 172 42810
rect 1666 42872 1700 42906
rect 138 42584 172 42618
rect 1666 42680 1700 42714
rect 138 42392 172 42426
rect 1666 42488 1700 42522
rect 138 42200 172 42234
rect 1666 42296 1700 42330
rect 138 42008 172 42042
rect 1666 42104 1700 42138
rect 138 41816 172 41850
rect 1666 41912 1700 41946
rect 138 41624 172 41658
rect 1666 41720 1700 41754
rect 138 41432 172 41466
rect 1666 41528 1700 41562
rect 138 41240 172 41274
rect 1666 41336 1700 41370
rect 138 41048 172 41082
rect 1666 41144 1700 41178
rect 138 40856 172 40890
rect 1666 40952 1700 40986
rect 138 40664 172 40698
rect 1666 40760 1700 40794
rect 138 40472 172 40506
rect 1666 40568 1700 40602
rect 138 40280 172 40314
rect 1666 40376 1700 40410
rect 138 40088 172 40122
rect 1666 40184 1700 40218
rect 138 39896 172 39930
rect 1666 39992 1700 40026
rect 138 39704 172 39738
rect 1666 39800 1700 39834
rect 138 39512 172 39546
rect 1666 39608 1700 39642
rect 138 39320 172 39354
rect 1666 39416 1700 39450
rect 138 39128 172 39162
rect 1666 39224 1700 39258
rect 138 38936 172 38970
rect 1666 39032 1700 39066
rect 138 38744 172 38778
rect 1666 38840 1700 38874
rect 138 38552 172 38586
rect 1666 38648 1700 38682
rect 138 38360 172 38394
rect 1666 38456 1700 38490
rect 138 38168 172 38202
rect 1666 38264 1700 38298
rect 138 37976 172 38010
rect 1666 38072 1700 38106
rect 138 37784 172 37818
rect 1666 37880 1700 37914
rect 138 37592 172 37626
rect 1666 37688 1700 37722
rect 138 37400 172 37434
rect 1666 37496 1700 37530
rect 138 37208 172 37242
rect 1666 37304 1700 37338
rect 138 37016 172 37050
rect 1666 37112 1700 37146
rect 138 36824 172 36858
rect 1666 36920 1700 36954
rect 138 36632 172 36666
rect 1666 36728 1700 36762
rect 138 36440 172 36474
rect 1666 36536 1700 36570
rect 138 36248 172 36282
rect 1666 36344 1700 36378
rect 138 36056 172 36090
rect 1666 36152 1700 36186
rect 138 35864 172 35898
rect 1666 35960 1700 35994
rect 138 35672 172 35706
rect 1666 35768 1700 35802
rect 138 35480 172 35514
rect 1666 35576 1700 35610
rect 138 35288 172 35322
rect 1666 35384 1700 35418
rect 138 35096 172 35130
rect 1666 35192 1700 35226
rect 138 34904 172 34938
rect 1666 35000 1700 35034
rect 138 34712 172 34746
rect 1666 34808 1700 34842
rect 138 34520 172 34554
rect 1666 34616 1700 34650
rect 138 34328 172 34362
rect 1666 34424 1700 34458
rect 138 34136 172 34170
rect 1666 34232 1700 34266
rect 138 33944 172 33978
rect 1666 34040 1700 34074
rect 138 33752 172 33786
rect 1666 33848 1700 33882
rect 138 33560 172 33594
rect 1666 33656 1700 33690
rect 138 33368 172 33402
rect 1666 33464 1700 33498
rect 138 33176 172 33210
rect 1666 33272 1700 33306
rect 138 32984 172 33018
rect 1666 33080 1700 33114
rect 138 32792 172 32826
rect 1666 32888 1700 32922
rect 138 32600 172 32634
rect 1666 32696 1700 32730
rect 138 32408 172 32442
rect 1666 32504 1700 32538
rect 138 32216 172 32250
rect 1666 32312 1700 32346
rect 138 32024 172 32058
rect 1666 32120 1700 32154
rect 138 31832 172 31866
rect 1666 31928 1700 31962
rect 138 31640 172 31674
rect 1666 31736 1700 31770
rect 138 31448 172 31482
rect 1666 31544 1700 31578
rect 138 31256 172 31290
rect 1666 31352 1700 31386
rect 138 31064 172 31098
rect 1666 31160 1700 31194
rect 138 30872 172 30906
rect 1666 30968 1700 31002
rect 138 30680 172 30714
rect 1666 30776 1700 30810
rect 138 30488 172 30522
rect 1666 30584 1700 30618
rect 138 30296 172 30330
rect 1666 30392 1700 30426
rect 138 30104 172 30138
rect 1666 30200 1700 30234
rect 138 29912 172 29946
rect 1666 30008 1700 30042
rect 138 29720 172 29754
rect 1666 29816 1700 29850
rect 138 29528 172 29562
rect 1666 29624 1700 29658
rect 138 29336 172 29370
rect 1666 29432 1700 29466
rect 138 29144 172 29178
rect 1666 29240 1700 29274
rect 138 28952 172 28986
rect 1666 29048 1700 29082
rect 138 28760 172 28794
rect 1666 28856 1700 28890
rect 138 28568 172 28602
rect 1666 28664 1700 28698
rect 138 28376 172 28410
rect 1666 28472 1700 28506
rect 138 28184 172 28218
rect 1666 28280 1700 28314
rect 138 27992 172 28026
rect 1666 28088 1700 28122
rect 138 27800 172 27834
rect 1666 27896 1700 27930
rect 138 27608 172 27642
rect 1666 27704 1700 27738
rect 138 27416 172 27450
rect 1666 27512 1700 27546
rect 138 27224 172 27258
rect 1666 27320 1700 27354
rect 138 27032 172 27066
rect 1666 27128 1700 27162
rect 138 26840 172 26874
rect 1666 26936 1700 26970
rect 138 26648 172 26682
rect 1666 26744 1700 26778
rect 138 26456 172 26490
rect 1666 26552 1700 26586
rect 138 26264 172 26298
rect 1666 26360 1700 26394
rect 138 26072 172 26106
rect 1666 26168 1700 26202
rect 138 25880 172 25914
rect 1666 25976 1700 26010
rect 138 25688 172 25722
rect 1666 25784 1700 25818
rect 138 25496 172 25530
rect 1666 25592 1700 25626
rect 138 25304 172 25338
rect 1666 25400 1700 25434
rect 138 25112 172 25146
rect 1666 25208 1700 25242
rect 138 24920 172 24954
rect 1666 25016 1700 25050
rect 138 24728 172 24762
rect 1666 24824 1700 24858
rect 138 24536 172 24570
rect 1666 24632 1700 24666
rect 138 24344 172 24378
rect 1666 24440 1700 24474
rect 138 24152 172 24186
rect 1666 24248 1700 24282
rect 138 23960 172 23994
rect 1666 24056 1700 24090
rect 138 23768 172 23802
rect 1666 23864 1700 23898
rect 138 23576 172 23610
rect 1666 23672 1700 23706
rect 138 23384 172 23418
rect 1666 23480 1700 23514
rect 138 23192 172 23226
rect 1666 23288 1700 23322
rect 1666 23096 1700 23130
rect 138 21622 172 21656
rect 138 21430 172 21464
rect 1666 21526 1700 21560
rect 138 21238 172 21272
rect 1666 21334 1700 21368
rect 138 21046 172 21080
rect 1666 21142 1700 21176
rect 138 20854 172 20888
rect 1666 20950 1700 20984
rect 138 20662 172 20696
rect 1666 20758 1700 20792
rect 138 20470 172 20504
rect 1666 20566 1700 20600
rect 138 20278 172 20312
rect 1666 20374 1700 20408
rect 138 20086 172 20120
rect 1666 20182 1700 20216
rect 138 19894 172 19928
rect 1666 19990 1700 20024
rect 138 19702 172 19736
rect 1666 19798 1700 19832
rect 138 19510 172 19544
rect 1666 19606 1700 19640
rect 138 19318 172 19352
rect 1666 19414 1700 19448
rect 138 19126 172 19160
rect 1666 19222 1700 19256
rect 138 18934 172 18968
rect 1666 19030 1700 19064
rect 138 18742 172 18776
rect 1666 18838 1700 18872
rect 138 18550 172 18584
rect 1666 18646 1700 18680
rect 138 18358 172 18392
rect 1666 18454 1700 18488
rect 138 18166 172 18200
rect 1666 18262 1700 18296
rect 138 17974 172 18008
rect 1666 18070 1700 18104
rect 138 17782 172 17816
rect 1666 17878 1700 17912
rect 138 17590 172 17624
rect 1666 17686 1700 17720
rect 138 17398 172 17432
rect 1666 17494 1700 17528
rect 138 17206 172 17240
rect 1666 17302 1700 17336
rect 138 17014 172 17048
rect 1666 17110 1700 17144
rect 138 16822 172 16856
rect 1666 16918 1700 16952
rect 138 16630 172 16664
rect 1666 16726 1700 16760
rect 138 16438 172 16472
rect 1666 16534 1700 16568
rect 138 16246 172 16280
rect 1666 16342 1700 16376
rect 138 16054 172 16088
rect 1666 16150 1700 16184
rect 138 15862 172 15896
rect 1666 15958 1700 15992
rect 138 15670 172 15704
rect 1666 15766 1700 15800
rect 138 15478 172 15512
rect 1666 15574 1700 15608
rect 138 15286 172 15320
rect 1666 15382 1700 15416
rect 138 15094 172 15128
rect 1666 15190 1700 15224
rect 138 14902 172 14936
rect 1666 14998 1700 15032
rect 138 14710 172 14744
rect 1666 14806 1700 14840
rect 138 14518 172 14552
rect 1666 14614 1700 14648
rect 138 14326 172 14360
rect 1666 14422 1700 14456
rect 138 14134 172 14168
rect 1666 14230 1700 14264
rect 138 13942 172 13976
rect 1666 14038 1700 14072
rect 138 13750 172 13784
rect 1666 13846 1700 13880
rect 138 13558 172 13592
rect 1666 13654 1700 13688
rect 138 13366 172 13400
rect 1666 13462 1700 13496
rect 138 13174 172 13208
rect 1666 13270 1700 13304
rect 138 12982 172 13016
rect 1666 13078 1700 13112
rect 138 12790 172 12824
rect 1666 12886 1700 12920
rect 138 12598 172 12632
rect 1666 12694 1700 12728
rect 138 12406 172 12440
rect 1666 12502 1700 12536
rect 138 12214 172 12248
rect 1666 12310 1700 12344
rect 138 12022 172 12056
rect 1666 12118 1700 12152
rect 138 11830 172 11864
rect 1666 11926 1700 11960
rect 138 11638 172 11672
rect 1666 11734 1700 11768
rect 138 11446 172 11480
rect 1666 11542 1700 11576
rect 138 11254 172 11288
rect 1666 11350 1700 11384
rect 138 11062 172 11096
rect 1666 11158 1700 11192
rect 138 10870 172 10904
rect 1666 10966 1700 11000
rect 138 10678 172 10712
rect 1666 10774 1700 10808
rect 138 10486 172 10520
rect 1666 10582 1700 10616
rect 138 10294 172 10328
rect 1666 10390 1700 10424
rect 138 10102 172 10136
rect 1666 10198 1700 10232
rect 138 9910 172 9944
rect 1666 10006 1700 10040
rect 138 9718 172 9752
rect 1666 9814 1700 9848
rect 138 9526 172 9560
rect 1666 9622 1700 9656
rect 138 9334 172 9368
rect 1666 9430 1700 9464
rect 138 9142 172 9176
rect 1666 9238 1700 9272
rect 138 8950 172 8984
rect 1666 9046 1700 9080
rect 138 8758 172 8792
rect 1666 8854 1700 8888
rect 138 8566 172 8600
rect 1666 8662 1700 8696
rect 138 8374 172 8408
rect 1666 8470 1700 8504
rect 138 8182 172 8216
rect 1666 8278 1700 8312
rect 138 7990 172 8024
rect 1666 8086 1700 8120
rect 138 7798 172 7832
rect 1666 7894 1700 7928
rect 138 7606 172 7640
rect 1666 7702 1700 7736
rect 138 7414 172 7448
rect 1666 7510 1700 7544
rect 138 7222 172 7256
rect 1666 7318 1700 7352
rect 138 7030 172 7064
rect 1666 7126 1700 7160
rect 138 6838 172 6872
rect 1666 6934 1700 6968
rect 138 6646 172 6680
rect 1666 6742 1700 6776
rect 138 6454 172 6488
rect 1666 6550 1700 6584
rect 138 6262 172 6296
rect 1666 6358 1700 6392
rect 138 6070 172 6104
rect 1666 6166 1700 6200
rect 138 5878 172 5912
rect 1666 5974 1700 6008
rect 138 5686 172 5720
rect 1666 5782 1700 5816
rect 138 5494 172 5528
rect 1666 5590 1700 5624
rect 138 5302 172 5336
rect 1666 5398 1700 5432
rect 138 5110 172 5144
rect 1666 5206 1700 5240
rect 138 4918 172 4952
rect 1666 5014 1700 5048
rect 138 4726 172 4760
rect 1666 4822 1700 4856
rect 138 4534 172 4568
rect 1666 4630 1700 4664
rect 138 4342 172 4376
rect 1666 4438 1700 4472
rect 138 4150 172 4184
rect 1666 4246 1700 4280
rect 138 3958 172 3992
rect 1666 4054 1700 4088
rect 138 3766 172 3800
rect 1666 3862 1700 3896
rect 138 3574 172 3608
rect 1666 3670 1700 3704
rect 138 3382 172 3416
rect 1666 3478 1700 3512
rect 138 3190 172 3224
rect 1666 3286 1700 3320
rect 138 2998 172 3032
rect 1666 3094 1700 3128
rect 138 2806 172 2840
rect 1666 2902 1700 2936
rect 138 2614 172 2648
rect 1666 2710 1700 2744
rect 138 2422 172 2456
rect 1666 2518 1700 2552
rect 138 2230 172 2264
rect 1666 2326 1700 2360
rect 138 2038 172 2072
rect 1666 2134 1700 2168
rect 138 1846 172 1880
rect 1666 1942 1700 1976
rect 138 1654 172 1688
rect 1666 1750 1700 1784
rect 138 1462 172 1496
rect 1666 1558 1700 1592
rect 138 1270 172 1304
rect 1666 1366 1700 1400
rect 138 1078 172 1112
rect 1666 1174 1700 1208
rect 138 886 172 920
rect 1666 982 1700 1016
rect 138 694 172 728
rect 1666 790 1700 824
rect 1666 598 1700 632
<< locali >>
rect 36 44282 132 44316
rect 1706 44282 1802 44316
rect 36 44220 70 44282
rect 1768 44220 1802 44282
rect 138 44154 172 44170
rect 215 44168 231 44202
rect 1607 44168 1623 44202
rect 138 44104 172 44120
rect 215 44072 231 44106
rect 1607 44072 1623 44106
rect 1666 44058 1700 44074
rect 138 43962 172 43978
rect 215 43976 231 44010
rect 1607 43976 1623 44010
rect 1666 44008 1700 44024
rect 138 43912 172 43928
rect 215 43880 231 43914
rect 1607 43880 1623 43914
rect 1666 43866 1700 43882
rect 138 43770 172 43786
rect 215 43784 231 43818
rect 1607 43784 1623 43818
rect 1666 43816 1700 43832
rect 138 43720 172 43736
rect 215 43688 231 43722
rect 1607 43688 1623 43722
rect 1666 43674 1700 43690
rect 138 43578 172 43594
rect 215 43592 231 43626
rect 1607 43592 1623 43626
rect 1666 43624 1700 43640
rect 138 43528 172 43544
rect 215 43496 231 43530
rect 1607 43496 1623 43530
rect 1666 43482 1700 43498
rect 138 43386 172 43402
rect 215 43400 231 43434
rect 1607 43400 1623 43434
rect 1666 43432 1700 43448
rect 138 43336 172 43352
rect 215 43304 231 43338
rect 1607 43304 1623 43338
rect 1666 43290 1700 43306
rect 138 43194 172 43210
rect 215 43208 231 43242
rect 1607 43208 1623 43242
rect 1666 43240 1700 43256
rect 138 43144 172 43160
rect 215 43112 231 43146
rect 1607 43112 1623 43146
rect 1666 43098 1700 43114
rect 138 43002 172 43018
rect 215 43016 231 43050
rect 1607 43016 1623 43050
rect 1666 43048 1700 43064
rect 138 42952 172 42968
rect 215 42920 231 42954
rect 1607 42920 1623 42954
rect 1666 42906 1700 42922
rect 138 42810 172 42826
rect 215 42824 231 42858
rect 1607 42824 1623 42858
rect 1666 42856 1700 42872
rect 138 42760 172 42776
rect 215 42728 231 42762
rect 1607 42728 1623 42762
rect 1666 42714 1700 42730
rect 138 42618 172 42634
rect 215 42632 231 42666
rect 1607 42632 1623 42666
rect 1666 42664 1700 42680
rect 138 42568 172 42584
rect 215 42536 231 42570
rect 1607 42536 1623 42570
rect 1666 42522 1700 42538
rect 138 42426 172 42442
rect 215 42440 231 42474
rect 1607 42440 1623 42474
rect 1666 42472 1700 42488
rect 138 42376 172 42392
rect 215 42344 231 42378
rect 1607 42344 1623 42378
rect 1666 42330 1700 42346
rect 138 42234 172 42250
rect 215 42248 231 42282
rect 1607 42248 1623 42282
rect 1666 42280 1700 42296
rect 138 42184 172 42200
rect 215 42152 231 42186
rect 1607 42152 1623 42186
rect 1666 42138 1700 42154
rect 138 42042 172 42058
rect 215 42056 231 42090
rect 1607 42056 1623 42090
rect 1666 42088 1700 42104
rect 138 41992 172 42008
rect 215 41960 231 41994
rect 1607 41960 1623 41994
rect 1666 41946 1700 41962
rect 138 41850 172 41866
rect 215 41864 231 41898
rect 1607 41864 1623 41898
rect 1666 41896 1700 41912
rect 138 41800 172 41816
rect 215 41768 231 41802
rect 1607 41768 1623 41802
rect 1666 41754 1700 41770
rect 138 41658 172 41674
rect 215 41672 231 41706
rect 1607 41672 1623 41706
rect 1666 41704 1700 41720
rect 138 41608 172 41624
rect 215 41576 231 41610
rect 1607 41576 1623 41610
rect 1666 41562 1700 41578
rect 138 41466 172 41482
rect 215 41480 231 41514
rect 1607 41480 1623 41514
rect 1666 41512 1700 41528
rect 138 41416 172 41432
rect 215 41384 231 41418
rect 1607 41384 1623 41418
rect 1666 41370 1700 41386
rect 138 41274 172 41290
rect 215 41288 231 41322
rect 1607 41288 1623 41322
rect 1666 41320 1700 41336
rect 138 41224 172 41240
rect 215 41192 231 41226
rect 1607 41192 1623 41226
rect 1666 41178 1700 41194
rect 138 41082 172 41098
rect 215 41096 231 41130
rect 1607 41096 1623 41130
rect 1666 41128 1700 41144
rect 138 41032 172 41048
rect 215 41000 231 41034
rect 1607 41000 1623 41034
rect 1666 40986 1700 41002
rect 138 40890 172 40906
rect 215 40904 231 40938
rect 1607 40904 1623 40938
rect 1666 40936 1700 40952
rect 138 40840 172 40856
rect 215 40808 231 40842
rect 1607 40808 1623 40842
rect 1666 40794 1700 40810
rect 138 40698 172 40714
rect 215 40712 231 40746
rect 1607 40712 1623 40746
rect 1666 40744 1700 40760
rect 138 40648 172 40664
rect 215 40616 231 40650
rect 1607 40616 1623 40650
rect 1666 40602 1700 40618
rect 138 40506 172 40522
rect 215 40520 231 40554
rect 1607 40520 1623 40554
rect 1666 40552 1700 40568
rect 138 40456 172 40472
rect 215 40424 231 40458
rect 1607 40424 1623 40458
rect 1666 40410 1700 40426
rect 138 40314 172 40330
rect 215 40328 231 40362
rect 1607 40328 1623 40362
rect 1666 40360 1700 40376
rect 138 40264 172 40280
rect 215 40232 231 40266
rect 1607 40232 1623 40266
rect 1666 40218 1700 40234
rect 138 40122 172 40138
rect 215 40136 231 40170
rect 1607 40136 1623 40170
rect 1666 40168 1700 40184
rect 138 40072 172 40088
rect 215 40040 231 40074
rect 1607 40040 1623 40074
rect 1666 40026 1700 40042
rect 138 39930 172 39946
rect 215 39944 231 39978
rect 1607 39944 1623 39978
rect 1666 39976 1700 39992
rect 138 39880 172 39896
rect 215 39848 231 39882
rect 1607 39848 1623 39882
rect 1666 39834 1700 39850
rect 138 39738 172 39754
rect 215 39752 231 39786
rect 1607 39752 1623 39786
rect 1666 39784 1700 39800
rect 138 39688 172 39704
rect 215 39656 231 39690
rect 1607 39656 1623 39690
rect 1666 39642 1700 39658
rect 138 39546 172 39562
rect 215 39560 231 39594
rect 1607 39560 1623 39594
rect 1666 39592 1700 39608
rect 138 39496 172 39512
rect 215 39464 231 39498
rect 1607 39464 1623 39498
rect 1666 39450 1700 39466
rect 138 39354 172 39370
rect 215 39368 231 39402
rect 1607 39368 1623 39402
rect 1666 39400 1700 39416
rect 138 39304 172 39320
rect 215 39272 231 39306
rect 1607 39272 1623 39306
rect 1666 39258 1700 39274
rect 138 39162 172 39178
rect 215 39176 231 39210
rect 1607 39176 1623 39210
rect 1666 39208 1700 39224
rect 138 39112 172 39128
rect 215 39080 231 39114
rect 1607 39080 1623 39114
rect 1666 39066 1700 39082
rect 138 38970 172 38986
rect 215 38984 231 39018
rect 1607 38984 1623 39018
rect 1666 39016 1700 39032
rect 138 38920 172 38936
rect 215 38888 231 38922
rect 1607 38888 1623 38922
rect 1666 38874 1700 38890
rect 138 38778 172 38794
rect 215 38792 231 38826
rect 1607 38792 1623 38826
rect 1666 38824 1700 38840
rect 138 38728 172 38744
rect 215 38696 231 38730
rect 1607 38696 1623 38730
rect 1666 38682 1700 38698
rect 138 38586 172 38602
rect 215 38600 231 38634
rect 1607 38600 1623 38634
rect 1666 38632 1700 38648
rect 138 38536 172 38552
rect 215 38504 231 38538
rect 1607 38504 1623 38538
rect 1666 38490 1700 38506
rect 138 38394 172 38410
rect 215 38408 231 38442
rect 1607 38408 1623 38442
rect 1666 38440 1700 38456
rect 138 38344 172 38360
rect 215 38312 231 38346
rect 1607 38312 1623 38346
rect 1666 38298 1700 38314
rect 138 38202 172 38218
rect 215 38216 231 38250
rect 1607 38216 1623 38250
rect 1666 38248 1700 38264
rect 138 38152 172 38168
rect 215 38120 231 38154
rect 1607 38120 1623 38154
rect 1666 38106 1700 38122
rect 138 38010 172 38026
rect 215 38024 231 38058
rect 1607 38024 1623 38058
rect 1666 38056 1700 38072
rect 138 37960 172 37976
rect 215 37928 231 37962
rect 1607 37928 1623 37962
rect 1666 37914 1700 37930
rect 138 37818 172 37834
rect 215 37832 231 37866
rect 1607 37832 1623 37866
rect 1666 37864 1700 37880
rect 138 37768 172 37784
rect 215 37736 231 37770
rect 1607 37736 1623 37770
rect 1666 37722 1700 37738
rect 138 37626 172 37642
rect 215 37640 231 37674
rect 1607 37640 1623 37674
rect 1666 37672 1700 37688
rect 138 37576 172 37592
rect 215 37544 231 37578
rect 1607 37544 1623 37578
rect 1666 37530 1700 37546
rect 138 37434 172 37450
rect 215 37448 231 37482
rect 1607 37448 1623 37482
rect 1666 37480 1700 37496
rect 138 37384 172 37400
rect 215 37352 231 37386
rect 1607 37352 1623 37386
rect 1666 37338 1700 37354
rect 138 37242 172 37258
rect 215 37256 231 37290
rect 1607 37256 1623 37290
rect 1666 37288 1700 37304
rect 138 37192 172 37208
rect 215 37160 231 37194
rect 1607 37160 1623 37194
rect 1666 37146 1700 37162
rect 138 37050 172 37066
rect 215 37064 231 37098
rect 1607 37064 1623 37098
rect 1666 37096 1700 37112
rect 138 37000 172 37016
rect 215 36968 231 37002
rect 1607 36968 1623 37002
rect 1666 36954 1700 36970
rect 138 36858 172 36874
rect 215 36872 231 36906
rect 1607 36872 1623 36906
rect 1666 36904 1700 36920
rect 138 36808 172 36824
rect 215 36776 231 36810
rect 1607 36776 1623 36810
rect 1666 36762 1700 36778
rect 138 36666 172 36682
rect 215 36680 231 36714
rect 1607 36680 1623 36714
rect 1666 36712 1700 36728
rect 138 36616 172 36632
rect 215 36584 231 36618
rect 1607 36584 1623 36618
rect 1666 36570 1700 36586
rect 138 36474 172 36490
rect 215 36488 231 36522
rect 1607 36488 1623 36522
rect 1666 36520 1700 36536
rect 138 36424 172 36440
rect 215 36392 231 36426
rect 1607 36392 1623 36426
rect 1666 36378 1700 36394
rect 138 36282 172 36298
rect 215 36296 231 36330
rect 1607 36296 1623 36330
rect 1666 36328 1700 36344
rect 138 36232 172 36248
rect 215 36200 231 36234
rect 1607 36200 1623 36234
rect 1666 36186 1700 36202
rect 138 36090 172 36106
rect 215 36104 231 36138
rect 1607 36104 1623 36138
rect 1666 36136 1700 36152
rect 138 36040 172 36056
rect 215 36008 231 36042
rect 1607 36008 1623 36042
rect 1666 35994 1700 36010
rect 138 35898 172 35914
rect 215 35912 231 35946
rect 1607 35912 1623 35946
rect 1666 35944 1700 35960
rect 138 35848 172 35864
rect 215 35816 231 35850
rect 1607 35816 1623 35850
rect 1666 35802 1700 35818
rect 138 35706 172 35722
rect 215 35720 231 35754
rect 1607 35720 1623 35754
rect 1666 35752 1700 35768
rect 138 35656 172 35672
rect 215 35624 231 35658
rect 1607 35624 1623 35658
rect 1666 35610 1700 35626
rect 138 35514 172 35530
rect 215 35528 231 35562
rect 1607 35528 1623 35562
rect 1666 35560 1700 35576
rect 138 35464 172 35480
rect 215 35432 231 35466
rect 1607 35432 1623 35466
rect 1666 35418 1700 35434
rect 138 35322 172 35338
rect 215 35336 231 35370
rect 1607 35336 1623 35370
rect 1666 35368 1700 35384
rect 138 35272 172 35288
rect 215 35240 231 35274
rect 1607 35240 1623 35274
rect 1666 35226 1700 35242
rect 138 35130 172 35146
rect 215 35144 231 35178
rect 1607 35144 1623 35178
rect 1666 35176 1700 35192
rect 138 35080 172 35096
rect 215 35048 231 35082
rect 1607 35048 1623 35082
rect 1666 35034 1700 35050
rect 138 34938 172 34954
rect 215 34952 231 34986
rect 1607 34952 1623 34986
rect 1666 34984 1700 35000
rect 138 34888 172 34904
rect 215 34856 231 34890
rect 1607 34856 1623 34890
rect 1666 34842 1700 34858
rect 138 34746 172 34762
rect 215 34760 231 34794
rect 1607 34760 1623 34794
rect 1666 34792 1700 34808
rect 138 34696 172 34712
rect 215 34664 231 34698
rect 1607 34664 1623 34698
rect 1666 34650 1700 34666
rect 138 34554 172 34570
rect 215 34568 231 34602
rect 1607 34568 1623 34602
rect 1666 34600 1700 34616
rect 138 34504 172 34520
rect 215 34472 231 34506
rect 1607 34472 1623 34506
rect 1666 34458 1700 34474
rect 138 34362 172 34378
rect 215 34376 231 34410
rect 1607 34376 1623 34410
rect 1666 34408 1700 34424
rect 138 34312 172 34328
rect 215 34280 231 34314
rect 1607 34280 1623 34314
rect 1666 34266 1700 34282
rect 138 34170 172 34186
rect 215 34184 231 34218
rect 1607 34184 1623 34218
rect 1666 34216 1700 34232
rect 138 34120 172 34136
rect 215 34088 231 34122
rect 1607 34088 1623 34122
rect 1666 34074 1700 34090
rect 138 33978 172 33994
rect 215 33992 231 34026
rect 1607 33992 1623 34026
rect 1666 34024 1700 34040
rect 138 33928 172 33944
rect 215 33896 231 33930
rect 1607 33896 1623 33930
rect 1666 33882 1700 33898
rect 138 33786 172 33802
rect 215 33800 231 33834
rect 1607 33800 1623 33834
rect 1666 33832 1700 33848
rect 138 33736 172 33752
rect 215 33704 231 33738
rect 1607 33704 1623 33738
rect 1666 33690 1700 33706
rect 138 33594 172 33610
rect 215 33608 231 33642
rect 1607 33608 1623 33642
rect 1666 33640 1700 33656
rect 138 33544 172 33560
rect 215 33512 231 33546
rect 1607 33512 1623 33546
rect 1666 33498 1700 33514
rect 138 33402 172 33418
rect 215 33416 231 33450
rect 1607 33416 1623 33450
rect 1666 33448 1700 33464
rect 138 33352 172 33368
rect 215 33320 231 33354
rect 1607 33320 1623 33354
rect 1666 33306 1700 33322
rect 138 33210 172 33226
rect 215 33224 231 33258
rect 1607 33224 1623 33258
rect 1666 33256 1700 33272
rect 138 33160 172 33176
rect 215 33128 231 33162
rect 1607 33128 1623 33162
rect 1666 33114 1700 33130
rect 138 33018 172 33034
rect 215 33032 231 33066
rect 1607 33032 1623 33066
rect 1666 33064 1700 33080
rect 138 32968 172 32984
rect 215 32936 231 32970
rect 1607 32936 1623 32970
rect 1666 32922 1700 32938
rect 138 32826 172 32842
rect 215 32840 231 32874
rect 1607 32840 1623 32874
rect 1666 32872 1700 32888
rect 138 32776 172 32792
rect 215 32744 231 32778
rect 1607 32744 1623 32778
rect 1666 32730 1700 32746
rect 138 32634 172 32650
rect 215 32648 231 32682
rect 1607 32648 1623 32682
rect 1666 32680 1700 32696
rect 138 32584 172 32600
rect 215 32552 231 32586
rect 1607 32552 1623 32586
rect 1666 32538 1700 32554
rect 138 32442 172 32458
rect 215 32456 231 32490
rect 1607 32456 1623 32490
rect 1666 32488 1700 32504
rect 138 32392 172 32408
rect 215 32360 231 32394
rect 1607 32360 1623 32394
rect 1666 32346 1700 32362
rect 138 32250 172 32266
rect 215 32264 231 32298
rect 1607 32264 1623 32298
rect 1666 32296 1700 32312
rect 138 32200 172 32216
rect 215 32168 231 32202
rect 1607 32168 1623 32202
rect 1666 32154 1700 32170
rect 138 32058 172 32074
rect 215 32072 231 32106
rect 1607 32072 1623 32106
rect 1666 32104 1700 32120
rect 138 32008 172 32024
rect 215 31976 231 32010
rect 1607 31976 1623 32010
rect 1666 31962 1700 31978
rect 138 31866 172 31882
rect 215 31880 231 31914
rect 1607 31880 1623 31914
rect 1666 31912 1700 31928
rect 138 31816 172 31832
rect 215 31784 231 31818
rect 1607 31784 1623 31818
rect 1666 31770 1700 31786
rect 138 31674 172 31690
rect 215 31688 231 31722
rect 1607 31688 1623 31722
rect 1666 31720 1700 31736
rect 138 31624 172 31640
rect 215 31592 231 31626
rect 1607 31592 1623 31626
rect 1666 31578 1700 31594
rect 138 31482 172 31498
rect 215 31496 231 31530
rect 1607 31496 1623 31530
rect 1666 31528 1700 31544
rect 138 31432 172 31448
rect 215 31400 231 31434
rect 1607 31400 1623 31434
rect 1666 31386 1700 31402
rect 138 31290 172 31306
rect 215 31304 231 31338
rect 1607 31304 1623 31338
rect 1666 31336 1700 31352
rect 138 31240 172 31256
rect 215 31208 231 31242
rect 1607 31208 1623 31242
rect 1666 31194 1700 31210
rect 138 31098 172 31114
rect 215 31112 231 31146
rect 1607 31112 1623 31146
rect 1666 31144 1700 31160
rect 138 31048 172 31064
rect 215 31016 231 31050
rect 1607 31016 1623 31050
rect 1666 31002 1700 31018
rect 138 30906 172 30922
rect 215 30920 231 30954
rect 1607 30920 1623 30954
rect 1666 30952 1700 30968
rect 138 30856 172 30872
rect 215 30824 231 30858
rect 1607 30824 1623 30858
rect 1666 30810 1700 30826
rect 138 30714 172 30730
rect 215 30728 231 30762
rect 1607 30728 1623 30762
rect 1666 30760 1700 30776
rect 138 30664 172 30680
rect 215 30632 231 30666
rect 1607 30632 1623 30666
rect 1666 30618 1700 30634
rect 138 30522 172 30538
rect 215 30536 231 30570
rect 1607 30536 1623 30570
rect 1666 30568 1700 30584
rect 138 30472 172 30488
rect 215 30440 231 30474
rect 1607 30440 1623 30474
rect 1666 30426 1700 30442
rect 138 30330 172 30346
rect 215 30344 231 30378
rect 1607 30344 1623 30378
rect 1666 30376 1700 30392
rect 138 30280 172 30296
rect 215 30248 231 30282
rect 1607 30248 1623 30282
rect 1666 30234 1700 30250
rect 138 30138 172 30154
rect 215 30152 231 30186
rect 1607 30152 1623 30186
rect 1666 30184 1700 30200
rect 138 30088 172 30104
rect 215 30056 231 30090
rect 1607 30056 1623 30090
rect 1666 30042 1700 30058
rect 138 29946 172 29962
rect 215 29960 231 29994
rect 1607 29960 1623 29994
rect 1666 29992 1700 30008
rect 138 29896 172 29912
rect 215 29864 231 29898
rect 1607 29864 1623 29898
rect 1666 29850 1700 29866
rect 138 29754 172 29770
rect 215 29768 231 29802
rect 1607 29768 1623 29802
rect 1666 29800 1700 29816
rect 138 29704 172 29720
rect 215 29672 231 29706
rect 1607 29672 1623 29706
rect 1666 29658 1700 29674
rect 138 29562 172 29578
rect 215 29576 231 29610
rect 1607 29576 1623 29610
rect 1666 29608 1700 29624
rect 138 29512 172 29528
rect 215 29480 231 29514
rect 1607 29480 1623 29514
rect 1666 29466 1700 29482
rect 138 29370 172 29386
rect 215 29384 231 29418
rect 1607 29384 1623 29418
rect 1666 29416 1700 29432
rect 138 29320 172 29336
rect 215 29288 231 29322
rect 1607 29288 1623 29322
rect 1666 29274 1700 29290
rect 138 29178 172 29194
rect 215 29192 231 29226
rect 1607 29192 1623 29226
rect 1666 29224 1700 29240
rect 138 29128 172 29144
rect 215 29096 231 29130
rect 1607 29096 1623 29130
rect 1666 29082 1700 29098
rect 138 28986 172 29002
rect 215 29000 231 29034
rect 1607 29000 1623 29034
rect 1666 29032 1700 29048
rect 138 28936 172 28952
rect 215 28904 231 28938
rect 1607 28904 1623 28938
rect 1666 28890 1700 28906
rect 138 28794 172 28810
rect 215 28808 231 28842
rect 1607 28808 1623 28842
rect 1666 28840 1700 28856
rect 138 28744 172 28760
rect 215 28712 231 28746
rect 1607 28712 1623 28746
rect 1666 28698 1700 28714
rect 138 28602 172 28618
rect 215 28616 231 28650
rect 1607 28616 1623 28650
rect 1666 28648 1700 28664
rect 138 28552 172 28568
rect 215 28520 231 28554
rect 1607 28520 1623 28554
rect 1666 28506 1700 28522
rect 138 28410 172 28426
rect 215 28424 231 28458
rect 1607 28424 1623 28458
rect 1666 28456 1700 28472
rect 138 28360 172 28376
rect 215 28328 231 28362
rect 1607 28328 1623 28362
rect 1666 28314 1700 28330
rect 138 28218 172 28234
rect 215 28232 231 28266
rect 1607 28232 1623 28266
rect 1666 28264 1700 28280
rect 138 28168 172 28184
rect 215 28136 231 28170
rect 1607 28136 1623 28170
rect 1666 28122 1700 28138
rect 138 28026 172 28042
rect 215 28040 231 28074
rect 1607 28040 1623 28074
rect 1666 28072 1700 28088
rect 138 27976 172 27992
rect 215 27944 231 27978
rect 1607 27944 1623 27978
rect 1666 27930 1700 27946
rect 138 27834 172 27850
rect 215 27848 231 27882
rect 1607 27848 1623 27882
rect 1666 27880 1700 27896
rect 138 27784 172 27800
rect 215 27752 231 27786
rect 1607 27752 1623 27786
rect 1666 27738 1700 27754
rect 138 27642 172 27658
rect 215 27656 231 27690
rect 1607 27656 1623 27690
rect 1666 27688 1700 27704
rect 138 27592 172 27608
rect 215 27560 231 27594
rect 1607 27560 1623 27594
rect 1666 27546 1700 27562
rect 138 27450 172 27466
rect 215 27464 231 27498
rect 1607 27464 1623 27498
rect 1666 27496 1700 27512
rect 138 27400 172 27416
rect 215 27368 231 27402
rect 1607 27368 1623 27402
rect 1666 27354 1700 27370
rect 138 27258 172 27274
rect 215 27272 231 27306
rect 1607 27272 1623 27306
rect 1666 27304 1700 27320
rect 138 27208 172 27224
rect 215 27176 231 27210
rect 1607 27176 1623 27210
rect 1666 27162 1700 27178
rect 138 27066 172 27082
rect 215 27080 231 27114
rect 1607 27080 1623 27114
rect 1666 27112 1700 27128
rect 138 27016 172 27032
rect 215 26984 231 27018
rect 1607 26984 1623 27018
rect 1666 26970 1700 26986
rect 138 26874 172 26890
rect 215 26888 231 26922
rect 1607 26888 1623 26922
rect 1666 26920 1700 26936
rect 138 26824 172 26840
rect 215 26792 231 26826
rect 1607 26792 1623 26826
rect 1666 26778 1700 26794
rect 138 26682 172 26698
rect 215 26696 231 26730
rect 1607 26696 1623 26730
rect 1666 26728 1700 26744
rect 138 26632 172 26648
rect 215 26600 231 26634
rect 1607 26600 1623 26634
rect 1666 26586 1700 26602
rect 138 26490 172 26506
rect 215 26504 231 26538
rect 1607 26504 1623 26538
rect 1666 26536 1700 26552
rect 138 26440 172 26456
rect 215 26408 231 26442
rect 1607 26408 1623 26442
rect 1666 26394 1700 26410
rect 138 26298 172 26314
rect 215 26312 231 26346
rect 1607 26312 1623 26346
rect 1666 26344 1700 26360
rect 138 26248 172 26264
rect 215 26216 231 26250
rect 1607 26216 1623 26250
rect 1666 26202 1700 26218
rect 138 26106 172 26122
rect 215 26120 231 26154
rect 1607 26120 1623 26154
rect 1666 26152 1700 26168
rect 138 26056 172 26072
rect 215 26024 231 26058
rect 1607 26024 1623 26058
rect 1666 26010 1700 26026
rect 138 25914 172 25930
rect 215 25928 231 25962
rect 1607 25928 1623 25962
rect 1666 25960 1700 25976
rect 138 25864 172 25880
rect 215 25832 231 25866
rect 1607 25832 1623 25866
rect 1666 25818 1700 25834
rect 138 25722 172 25738
rect 215 25736 231 25770
rect 1607 25736 1623 25770
rect 1666 25768 1700 25784
rect 138 25672 172 25688
rect 215 25640 231 25674
rect 1607 25640 1623 25674
rect 1666 25626 1700 25642
rect 138 25530 172 25546
rect 215 25544 231 25578
rect 1607 25544 1623 25578
rect 1666 25576 1700 25592
rect 138 25480 172 25496
rect 215 25448 231 25482
rect 1607 25448 1623 25482
rect 1666 25434 1700 25450
rect 138 25338 172 25354
rect 215 25352 231 25386
rect 1607 25352 1623 25386
rect 1666 25384 1700 25400
rect 138 25288 172 25304
rect 215 25256 231 25290
rect 1607 25256 1623 25290
rect 1666 25242 1700 25258
rect 138 25146 172 25162
rect 215 25160 231 25194
rect 1607 25160 1623 25194
rect 1666 25192 1700 25208
rect 138 25096 172 25112
rect 215 25064 231 25098
rect 1607 25064 1623 25098
rect 1666 25050 1700 25066
rect 138 24954 172 24970
rect 215 24968 231 25002
rect 1607 24968 1623 25002
rect 1666 25000 1700 25016
rect 138 24904 172 24920
rect 215 24872 231 24906
rect 1607 24872 1623 24906
rect 1666 24858 1700 24874
rect 138 24762 172 24778
rect 215 24776 231 24810
rect 1607 24776 1623 24810
rect 1666 24808 1700 24824
rect 138 24712 172 24728
rect 215 24680 231 24714
rect 1607 24680 1623 24714
rect 1666 24666 1700 24682
rect 138 24570 172 24586
rect 215 24584 231 24618
rect 1607 24584 1623 24618
rect 1666 24616 1700 24632
rect 138 24520 172 24536
rect 215 24488 231 24522
rect 1607 24488 1623 24522
rect 1666 24474 1700 24490
rect 138 24378 172 24394
rect 215 24392 231 24426
rect 1607 24392 1623 24426
rect 1666 24424 1700 24440
rect 138 24328 172 24344
rect 215 24296 231 24330
rect 1607 24296 1623 24330
rect 1666 24282 1700 24298
rect 138 24186 172 24202
rect 215 24200 231 24234
rect 1607 24200 1623 24234
rect 1666 24232 1700 24248
rect 138 24136 172 24152
rect 215 24104 231 24138
rect 1607 24104 1623 24138
rect 1666 24090 1700 24106
rect 138 23994 172 24010
rect 215 24008 231 24042
rect 1607 24008 1623 24042
rect 1666 24040 1700 24056
rect 138 23944 172 23960
rect 215 23912 231 23946
rect 1607 23912 1623 23946
rect 1666 23898 1700 23914
rect 138 23802 172 23818
rect 215 23816 231 23850
rect 1607 23816 1623 23850
rect 1666 23848 1700 23864
rect 138 23752 172 23768
rect 215 23720 231 23754
rect 1607 23720 1623 23754
rect 1666 23706 1700 23722
rect 138 23610 172 23626
rect 215 23624 231 23658
rect 1607 23624 1623 23658
rect 1666 23656 1700 23672
rect 138 23560 172 23576
rect 215 23528 231 23562
rect 1607 23528 1623 23562
rect 1666 23514 1700 23530
rect 138 23418 172 23434
rect 215 23432 231 23466
rect 1607 23432 1623 23466
rect 1666 23464 1700 23480
rect 138 23368 172 23384
rect 215 23336 231 23370
rect 1607 23336 1623 23370
rect 1666 23322 1700 23338
rect 138 23226 172 23242
rect 215 23240 231 23274
rect 1607 23240 1623 23274
rect 1666 23272 1700 23288
rect 138 23176 172 23192
rect 215 23144 231 23178
rect 1607 23144 1623 23178
rect 1666 23130 1700 23146
rect 215 23048 231 23082
rect 1607 23048 1623 23082
rect 1666 23080 1700 23096
rect 36 22968 70 23030
rect 1768 22968 1802 23030
rect 36 22934 132 22968
rect 1706 22934 1802 22968
rect 36 22768 1802 22934
rect 36 21986 340 22768
rect 870 21986 1802 22768
rect 36 21818 1802 21986
rect 36 21784 132 21818
rect 1706 21784 1802 21818
rect 36 21722 70 21784
rect 1768 21722 1802 21784
rect 138 21656 172 21672
rect 215 21670 231 21704
rect 1607 21670 1623 21704
rect 138 21606 172 21622
rect 215 21574 231 21608
rect 1607 21574 1623 21608
rect 1666 21560 1700 21576
rect 138 21464 172 21480
rect 215 21478 231 21512
rect 1607 21478 1623 21512
rect 1666 21510 1700 21526
rect 138 21414 172 21430
rect 215 21382 231 21416
rect 1607 21382 1623 21416
rect 1666 21368 1700 21384
rect 138 21272 172 21288
rect 215 21286 231 21320
rect 1607 21286 1623 21320
rect 1666 21318 1700 21334
rect 138 21222 172 21238
rect 215 21190 231 21224
rect 1607 21190 1623 21224
rect 1666 21176 1700 21192
rect 138 21080 172 21096
rect 215 21094 231 21128
rect 1607 21094 1623 21128
rect 1666 21126 1700 21142
rect 138 21030 172 21046
rect 215 20998 231 21032
rect 1607 20998 1623 21032
rect 1666 20984 1700 21000
rect 138 20888 172 20904
rect 215 20902 231 20936
rect 1607 20902 1623 20936
rect 1666 20934 1700 20950
rect 138 20838 172 20854
rect 215 20806 231 20840
rect 1607 20806 1623 20840
rect 1666 20792 1700 20808
rect 138 20696 172 20712
rect 215 20710 231 20744
rect 1607 20710 1623 20744
rect 1666 20742 1700 20758
rect 138 20646 172 20662
rect 215 20614 231 20648
rect 1607 20614 1623 20648
rect 1666 20600 1700 20616
rect 138 20504 172 20520
rect 215 20518 231 20552
rect 1607 20518 1623 20552
rect 1666 20550 1700 20566
rect 138 20454 172 20470
rect 215 20422 231 20456
rect 1607 20422 1623 20456
rect 1666 20408 1700 20424
rect 138 20312 172 20328
rect 215 20326 231 20360
rect 1607 20326 1623 20360
rect 1666 20358 1700 20374
rect 138 20262 172 20278
rect 215 20230 231 20264
rect 1607 20230 1623 20264
rect 1666 20216 1700 20232
rect 138 20120 172 20136
rect 215 20134 231 20168
rect 1607 20134 1623 20168
rect 1666 20166 1700 20182
rect 138 20070 172 20086
rect 215 20038 231 20072
rect 1607 20038 1623 20072
rect 1666 20024 1700 20040
rect 138 19928 172 19944
rect 215 19942 231 19976
rect 1607 19942 1623 19976
rect 1666 19974 1700 19990
rect 138 19878 172 19894
rect 215 19846 231 19880
rect 1607 19846 1623 19880
rect 1666 19832 1700 19848
rect 138 19736 172 19752
rect 215 19750 231 19784
rect 1607 19750 1623 19784
rect 1666 19782 1700 19798
rect 138 19686 172 19702
rect 215 19654 231 19688
rect 1607 19654 1623 19688
rect 1666 19640 1700 19656
rect 138 19544 172 19560
rect 215 19558 231 19592
rect 1607 19558 1623 19592
rect 1666 19590 1700 19606
rect 138 19494 172 19510
rect 215 19462 231 19496
rect 1607 19462 1623 19496
rect 1666 19448 1700 19464
rect 138 19352 172 19368
rect 215 19366 231 19400
rect 1607 19366 1623 19400
rect 1666 19398 1700 19414
rect 138 19302 172 19318
rect 215 19270 231 19304
rect 1607 19270 1623 19304
rect 1666 19256 1700 19272
rect 138 19160 172 19176
rect 215 19174 231 19208
rect 1607 19174 1623 19208
rect 1666 19206 1700 19222
rect 138 19110 172 19126
rect 215 19078 231 19112
rect 1607 19078 1623 19112
rect 1666 19064 1700 19080
rect 138 18968 172 18984
rect 215 18982 231 19016
rect 1607 18982 1623 19016
rect 1666 19014 1700 19030
rect 138 18918 172 18934
rect 215 18886 231 18920
rect 1607 18886 1623 18920
rect 1666 18872 1700 18888
rect 138 18776 172 18792
rect 215 18790 231 18824
rect 1607 18790 1623 18824
rect 1666 18822 1700 18838
rect 138 18726 172 18742
rect 215 18694 231 18728
rect 1607 18694 1623 18728
rect 1666 18680 1700 18696
rect 138 18584 172 18600
rect 215 18598 231 18632
rect 1607 18598 1623 18632
rect 1666 18630 1700 18646
rect 138 18534 172 18550
rect 215 18502 231 18536
rect 1607 18502 1623 18536
rect 1666 18488 1700 18504
rect 138 18392 172 18408
rect 215 18406 231 18440
rect 1607 18406 1623 18440
rect 1666 18438 1700 18454
rect 138 18342 172 18358
rect 215 18310 231 18344
rect 1607 18310 1623 18344
rect 1666 18296 1700 18312
rect 138 18200 172 18216
rect 215 18214 231 18248
rect 1607 18214 1623 18248
rect 1666 18246 1700 18262
rect 138 18150 172 18166
rect 215 18118 231 18152
rect 1607 18118 1623 18152
rect 1666 18104 1700 18120
rect 138 18008 172 18024
rect 215 18022 231 18056
rect 1607 18022 1623 18056
rect 1666 18054 1700 18070
rect 138 17958 172 17974
rect 215 17926 231 17960
rect 1607 17926 1623 17960
rect 1666 17912 1700 17928
rect 138 17816 172 17832
rect 215 17830 231 17864
rect 1607 17830 1623 17864
rect 1666 17862 1700 17878
rect 138 17766 172 17782
rect 215 17734 231 17768
rect 1607 17734 1623 17768
rect 1666 17720 1700 17736
rect 138 17624 172 17640
rect 215 17638 231 17672
rect 1607 17638 1623 17672
rect 1666 17670 1700 17686
rect 138 17574 172 17590
rect 215 17542 231 17576
rect 1607 17542 1623 17576
rect 1666 17528 1700 17544
rect 138 17432 172 17448
rect 215 17446 231 17480
rect 1607 17446 1623 17480
rect 1666 17478 1700 17494
rect 138 17382 172 17398
rect 215 17350 231 17384
rect 1607 17350 1623 17384
rect 1666 17336 1700 17352
rect 138 17240 172 17256
rect 215 17254 231 17288
rect 1607 17254 1623 17288
rect 1666 17286 1700 17302
rect 138 17190 172 17206
rect 215 17158 231 17192
rect 1607 17158 1623 17192
rect 1666 17144 1700 17160
rect 138 17048 172 17064
rect 215 17062 231 17096
rect 1607 17062 1623 17096
rect 1666 17094 1700 17110
rect 138 16998 172 17014
rect 215 16966 231 17000
rect 1607 16966 1623 17000
rect 1666 16952 1700 16968
rect 138 16856 172 16872
rect 215 16870 231 16904
rect 1607 16870 1623 16904
rect 1666 16902 1700 16918
rect 138 16806 172 16822
rect 215 16774 231 16808
rect 1607 16774 1623 16808
rect 1666 16760 1700 16776
rect 138 16664 172 16680
rect 215 16678 231 16712
rect 1607 16678 1623 16712
rect 1666 16710 1700 16726
rect 138 16614 172 16630
rect 215 16582 231 16616
rect 1607 16582 1623 16616
rect 1666 16568 1700 16584
rect 138 16472 172 16488
rect 215 16486 231 16520
rect 1607 16486 1623 16520
rect 1666 16518 1700 16534
rect 138 16422 172 16438
rect 215 16390 231 16424
rect 1607 16390 1623 16424
rect 1666 16376 1700 16392
rect 138 16280 172 16296
rect 215 16294 231 16328
rect 1607 16294 1623 16328
rect 1666 16326 1700 16342
rect 138 16230 172 16246
rect 215 16198 231 16232
rect 1607 16198 1623 16232
rect 1666 16184 1700 16200
rect 138 16088 172 16104
rect 215 16102 231 16136
rect 1607 16102 1623 16136
rect 1666 16134 1700 16150
rect 138 16038 172 16054
rect 215 16006 231 16040
rect 1607 16006 1623 16040
rect 1666 15992 1700 16008
rect 138 15896 172 15912
rect 215 15910 231 15944
rect 1607 15910 1623 15944
rect 1666 15942 1700 15958
rect 138 15846 172 15862
rect 215 15814 231 15848
rect 1607 15814 1623 15848
rect 1666 15800 1700 15816
rect 138 15704 172 15720
rect 215 15718 231 15752
rect 1607 15718 1623 15752
rect 1666 15750 1700 15766
rect 138 15654 172 15670
rect 215 15622 231 15656
rect 1607 15622 1623 15656
rect 1666 15608 1700 15624
rect 138 15512 172 15528
rect 215 15526 231 15560
rect 1607 15526 1623 15560
rect 1666 15558 1700 15574
rect 138 15462 172 15478
rect 215 15430 231 15464
rect 1607 15430 1623 15464
rect 1666 15416 1700 15432
rect 138 15320 172 15336
rect 215 15334 231 15368
rect 1607 15334 1623 15368
rect 1666 15366 1700 15382
rect 138 15270 172 15286
rect 215 15238 231 15272
rect 1607 15238 1623 15272
rect 1666 15224 1700 15240
rect 138 15128 172 15144
rect 215 15142 231 15176
rect 1607 15142 1623 15176
rect 1666 15174 1700 15190
rect 138 15078 172 15094
rect 215 15046 231 15080
rect 1607 15046 1623 15080
rect 1666 15032 1700 15048
rect 138 14936 172 14952
rect 215 14950 231 14984
rect 1607 14950 1623 14984
rect 1666 14982 1700 14998
rect 138 14886 172 14902
rect 215 14854 231 14888
rect 1607 14854 1623 14888
rect 1666 14840 1700 14856
rect 138 14744 172 14760
rect 215 14758 231 14792
rect 1607 14758 1623 14792
rect 1666 14790 1700 14806
rect 138 14694 172 14710
rect 215 14662 231 14696
rect 1607 14662 1623 14696
rect 1666 14648 1700 14664
rect 138 14552 172 14568
rect 215 14566 231 14600
rect 1607 14566 1623 14600
rect 1666 14598 1700 14614
rect 138 14502 172 14518
rect 215 14470 231 14504
rect 1607 14470 1623 14504
rect 1666 14456 1700 14472
rect 138 14360 172 14376
rect 215 14374 231 14408
rect 1607 14374 1623 14408
rect 1666 14406 1700 14422
rect 138 14310 172 14326
rect 215 14278 231 14312
rect 1607 14278 1623 14312
rect 1666 14264 1700 14280
rect 138 14168 172 14184
rect 215 14182 231 14216
rect 1607 14182 1623 14216
rect 1666 14214 1700 14230
rect 138 14118 172 14134
rect 215 14086 231 14120
rect 1607 14086 1623 14120
rect 1666 14072 1700 14088
rect 138 13976 172 13992
rect 215 13990 231 14024
rect 1607 13990 1623 14024
rect 1666 14022 1700 14038
rect 138 13926 172 13942
rect 215 13894 231 13928
rect 1607 13894 1623 13928
rect 1666 13880 1700 13896
rect 138 13784 172 13800
rect 215 13798 231 13832
rect 1607 13798 1623 13832
rect 1666 13830 1700 13846
rect 138 13734 172 13750
rect 215 13702 231 13736
rect 1607 13702 1623 13736
rect 1666 13688 1700 13704
rect 138 13592 172 13608
rect 215 13606 231 13640
rect 1607 13606 1623 13640
rect 1666 13638 1700 13654
rect 138 13542 172 13558
rect 215 13510 231 13544
rect 1607 13510 1623 13544
rect 1666 13496 1700 13512
rect 138 13400 172 13416
rect 215 13414 231 13448
rect 1607 13414 1623 13448
rect 1666 13446 1700 13462
rect 138 13350 172 13366
rect 215 13318 231 13352
rect 1607 13318 1623 13352
rect 1666 13304 1700 13320
rect 138 13208 172 13224
rect 215 13222 231 13256
rect 1607 13222 1623 13256
rect 1666 13254 1700 13270
rect 138 13158 172 13174
rect 215 13126 231 13160
rect 1607 13126 1623 13160
rect 1666 13112 1700 13128
rect 138 13016 172 13032
rect 215 13030 231 13064
rect 1607 13030 1623 13064
rect 1666 13062 1700 13078
rect 138 12966 172 12982
rect 215 12934 231 12968
rect 1607 12934 1623 12968
rect 1666 12920 1700 12936
rect 138 12824 172 12840
rect 215 12838 231 12872
rect 1607 12838 1623 12872
rect 1666 12870 1700 12886
rect 138 12774 172 12790
rect 215 12742 231 12776
rect 1607 12742 1623 12776
rect 1666 12728 1700 12744
rect 138 12632 172 12648
rect 215 12646 231 12680
rect 1607 12646 1623 12680
rect 1666 12678 1700 12694
rect 138 12582 172 12598
rect 215 12550 231 12584
rect 1607 12550 1623 12584
rect 1666 12536 1700 12552
rect 138 12440 172 12456
rect 215 12454 231 12488
rect 1607 12454 1623 12488
rect 1666 12486 1700 12502
rect 138 12390 172 12406
rect 215 12358 231 12392
rect 1607 12358 1623 12392
rect 1666 12344 1700 12360
rect 138 12248 172 12264
rect 215 12262 231 12296
rect 1607 12262 1623 12296
rect 1666 12294 1700 12310
rect 138 12198 172 12214
rect 215 12166 231 12200
rect 1607 12166 1623 12200
rect 1666 12152 1700 12168
rect 138 12056 172 12072
rect 215 12070 231 12104
rect 1607 12070 1623 12104
rect 1666 12102 1700 12118
rect 138 12006 172 12022
rect 215 11974 231 12008
rect 1607 11974 1623 12008
rect 1666 11960 1700 11976
rect 138 11864 172 11880
rect 215 11878 231 11912
rect 1607 11878 1623 11912
rect 1666 11910 1700 11926
rect 138 11814 172 11830
rect 215 11782 231 11816
rect 1607 11782 1623 11816
rect 1666 11768 1700 11784
rect 138 11672 172 11688
rect 215 11686 231 11720
rect 1607 11686 1623 11720
rect 1666 11718 1700 11734
rect 138 11622 172 11638
rect 215 11590 231 11624
rect 1607 11590 1623 11624
rect 1666 11576 1700 11592
rect 138 11480 172 11496
rect 215 11494 231 11528
rect 1607 11494 1623 11528
rect 1666 11526 1700 11542
rect 138 11430 172 11446
rect 215 11398 231 11432
rect 1607 11398 1623 11432
rect 1666 11384 1700 11400
rect 138 11288 172 11304
rect 215 11302 231 11336
rect 1607 11302 1623 11336
rect 1666 11334 1700 11350
rect 138 11238 172 11254
rect 215 11206 231 11240
rect 1607 11206 1623 11240
rect 1666 11192 1700 11208
rect 138 11096 172 11112
rect 215 11110 231 11144
rect 1607 11110 1623 11144
rect 1666 11142 1700 11158
rect 138 11046 172 11062
rect 215 11014 231 11048
rect 1607 11014 1623 11048
rect 1666 11000 1700 11016
rect 138 10904 172 10920
rect 215 10918 231 10952
rect 1607 10918 1623 10952
rect 1666 10950 1700 10966
rect 138 10854 172 10870
rect 215 10822 231 10856
rect 1607 10822 1623 10856
rect 1666 10808 1700 10824
rect 138 10712 172 10728
rect 215 10726 231 10760
rect 1607 10726 1623 10760
rect 1666 10758 1700 10774
rect 138 10662 172 10678
rect 215 10630 231 10664
rect 1607 10630 1623 10664
rect 1666 10616 1700 10632
rect 138 10520 172 10536
rect 215 10534 231 10568
rect 1607 10534 1623 10568
rect 1666 10566 1700 10582
rect 138 10470 172 10486
rect 215 10438 231 10472
rect 1607 10438 1623 10472
rect 1666 10424 1700 10440
rect 138 10328 172 10344
rect 215 10342 231 10376
rect 1607 10342 1623 10376
rect 1666 10374 1700 10390
rect 138 10278 172 10294
rect 215 10246 231 10280
rect 1607 10246 1623 10280
rect 1666 10232 1700 10248
rect 138 10136 172 10152
rect 215 10150 231 10184
rect 1607 10150 1623 10184
rect 1666 10182 1700 10198
rect 138 10086 172 10102
rect 215 10054 231 10088
rect 1607 10054 1623 10088
rect 1666 10040 1700 10056
rect 138 9944 172 9960
rect 215 9958 231 9992
rect 1607 9958 1623 9992
rect 1666 9990 1700 10006
rect 138 9894 172 9910
rect 215 9862 231 9896
rect 1607 9862 1623 9896
rect 1666 9848 1700 9864
rect 138 9752 172 9768
rect 215 9766 231 9800
rect 1607 9766 1623 9800
rect 1666 9798 1700 9814
rect 138 9702 172 9718
rect 215 9670 231 9704
rect 1607 9670 1623 9704
rect 1666 9656 1700 9672
rect 138 9560 172 9576
rect 215 9574 231 9608
rect 1607 9574 1623 9608
rect 1666 9606 1700 9622
rect 138 9510 172 9526
rect 215 9478 231 9512
rect 1607 9478 1623 9512
rect 1666 9464 1700 9480
rect 138 9368 172 9384
rect 215 9382 231 9416
rect 1607 9382 1623 9416
rect 1666 9414 1700 9430
rect 138 9318 172 9334
rect 215 9286 231 9320
rect 1607 9286 1623 9320
rect 1666 9272 1700 9288
rect 138 9176 172 9192
rect 215 9190 231 9224
rect 1607 9190 1623 9224
rect 1666 9222 1700 9238
rect 138 9126 172 9142
rect 215 9094 231 9128
rect 1607 9094 1623 9128
rect 1666 9080 1700 9096
rect 138 8984 172 9000
rect 215 8998 231 9032
rect 1607 8998 1623 9032
rect 1666 9030 1700 9046
rect 138 8934 172 8950
rect 215 8902 231 8936
rect 1607 8902 1623 8936
rect 1666 8888 1700 8904
rect 138 8792 172 8808
rect 215 8806 231 8840
rect 1607 8806 1623 8840
rect 1666 8838 1700 8854
rect 138 8742 172 8758
rect 215 8710 231 8744
rect 1607 8710 1623 8744
rect 1666 8696 1700 8712
rect 138 8600 172 8616
rect 215 8614 231 8648
rect 1607 8614 1623 8648
rect 1666 8646 1700 8662
rect 138 8550 172 8566
rect 215 8518 231 8552
rect 1607 8518 1623 8552
rect 1666 8504 1700 8520
rect 138 8408 172 8424
rect 215 8422 231 8456
rect 1607 8422 1623 8456
rect 1666 8454 1700 8470
rect 138 8358 172 8374
rect 215 8326 231 8360
rect 1607 8326 1623 8360
rect 1666 8312 1700 8328
rect 138 8216 172 8232
rect 215 8230 231 8264
rect 1607 8230 1623 8264
rect 1666 8262 1700 8278
rect 138 8166 172 8182
rect 215 8134 231 8168
rect 1607 8134 1623 8168
rect 1666 8120 1700 8136
rect 138 8024 172 8040
rect 215 8038 231 8072
rect 1607 8038 1623 8072
rect 1666 8070 1700 8086
rect 138 7974 172 7990
rect 215 7942 231 7976
rect 1607 7942 1623 7976
rect 1666 7928 1700 7944
rect 138 7832 172 7848
rect 215 7846 231 7880
rect 1607 7846 1623 7880
rect 1666 7878 1700 7894
rect 138 7782 172 7798
rect 215 7750 231 7784
rect 1607 7750 1623 7784
rect 1666 7736 1700 7752
rect 138 7640 172 7656
rect 215 7654 231 7688
rect 1607 7654 1623 7688
rect 1666 7686 1700 7702
rect 138 7590 172 7606
rect 215 7558 231 7592
rect 1607 7558 1623 7592
rect 1666 7544 1700 7560
rect 138 7448 172 7464
rect 215 7462 231 7496
rect 1607 7462 1623 7496
rect 1666 7494 1700 7510
rect 138 7398 172 7414
rect 215 7366 231 7400
rect 1607 7366 1623 7400
rect 1666 7352 1700 7368
rect 138 7256 172 7272
rect 215 7270 231 7304
rect 1607 7270 1623 7304
rect 1666 7302 1700 7318
rect 138 7206 172 7222
rect 215 7174 231 7208
rect 1607 7174 1623 7208
rect 1666 7160 1700 7176
rect 138 7064 172 7080
rect 215 7078 231 7112
rect 1607 7078 1623 7112
rect 1666 7110 1700 7126
rect 138 7014 172 7030
rect 215 6982 231 7016
rect 1607 6982 1623 7016
rect 1666 6968 1700 6984
rect 138 6872 172 6888
rect 215 6886 231 6920
rect 1607 6886 1623 6920
rect 1666 6918 1700 6934
rect 138 6822 172 6838
rect 215 6790 231 6824
rect 1607 6790 1623 6824
rect 1666 6776 1700 6792
rect 138 6680 172 6696
rect 215 6694 231 6728
rect 1607 6694 1623 6728
rect 1666 6726 1700 6742
rect 138 6630 172 6646
rect 215 6598 231 6632
rect 1607 6598 1623 6632
rect 1666 6584 1700 6600
rect 138 6488 172 6504
rect 215 6502 231 6536
rect 1607 6502 1623 6536
rect 1666 6534 1700 6550
rect 138 6438 172 6454
rect 215 6406 231 6440
rect 1607 6406 1623 6440
rect 1666 6392 1700 6408
rect 138 6296 172 6312
rect 215 6310 231 6344
rect 1607 6310 1623 6344
rect 1666 6342 1700 6358
rect 138 6246 172 6262
rect 215 6214 231 6248
rect 1607 6214 1623 6248
rect 1666 6200 1700 6216
rect 138 6104 172 6120
rect 215 6118 231 6152
rect 1607 6118 1623 6152
rect 1666 6150 1700 6166
rect 138 6054 172 6070
rect 215 6022 231 6056
rect 1607 6022 1623 6056
rect 1666 6008 1700 6024
rect 138 5912 172 5928
rect 215 5926 231 5960
rect 1607 5926 1623 5960
rect 1666 5958 1700 5974
rect 138 5862 172 5878
rect 215 5830 231 5864
rect 1607 5830 1623 5864
rect 1666 5816 1700 5832
rect 138 5720 172 5736
rect 215 5734 231 5768
rect 1607 5734 1623 5768
rect 1666 5766 1700 5782
rect 138 5670 172 5686
rect 215 5638 231 5672
rect 1607 5638 1623 5672
rect 1666 5624 1700 5640
rect 138 5528 172 5544
rect 215 5542 231 5576
rect 1607 5542 1623 5576
rect 1666 5574 1700 5590
rect 138 5478 172 5494
rect 215 5446 231 5480
rect 1607 5446 1623 5480
rect 1666 5432 1700 5448
rect 138 5336 172 5352
rect 215 5350 231 5384
rect 1607 5350 1623 5384
rect 1666 5382 1700 5398
rect 138 5286 172 5302
rect 215 5254 231 5288
rect 1607 5254 1623 5288
rect 1666 5240 1700 5256
rect 138 5144 172 5160
rect 215 5158 231 5192
rect 1607 5158 1623 5192
rect 1666 5190 1700 5206
rect 138 5094 172 5110
rect 215 5062 231 5096
rect 1607 5062 1623 5096
rect 1666 5048 1700 5064
rect 138 4952 172 4968
rect 215 4966 231 5000
rect 1607 4966 1623 5000
rect 1666 4998 1700 5014
rect 138 4902 172 4918
rect 215 4870 231 4904
rect 1607 4870 1623 4904
rect 1666 4856 1700 4872
rect 138 4760 172 4776
rect 215 4774 231 4808
rect 1607 4774 1623 4808
rect 1666 4806 1700 4822
rect 138 4710 172 4726
rect 215 4678 231 4712
rect 1607 4678 1623 4712
rect 1666 4664 1700 4680
rect 138 4568 172 4584
rect 215 4582 231 4616
rect 1607 4582 1623 4616
rect 1666 4614 1700 4630
rect 138 4518 172 4534
rect 215 4486 231 4520
rect 1607 4486 1623 4520
rect 1666 4472 1700 4488
rect 138 4376 172 4392
rect 215 4390 231 4424
rect 1607 4390 1623 4424
rect 1666 4422 1700 4438
rect 138 4326 172 4342
rect 215 4294 231 4328
rect 1607 4294 1623 4328
rect 1666 4280 1700 4296
rect 138 4184 172 4200
rect 215 4198 231 4232
rect 1607 4198 1623 4232
rect 1666 4230 1700 4246
rect 138 4134 172 4150
rect 215 4102 231 4136
rect 1607 4102 1623 4136
rect 1666 4088 1700 4104
rect 138 3992 172 4008
rect 215 4006 231 4040
rect 1607 4006 1623 4040
rect 1666 4038 1700 4054
rect 138 3942 172 3958
rect 215 3910 231 3944
rect 1607 3910 1623 3944
rect 1666 3896 1700 3912
rect 138 3800 172 3816
rect 215 3814 231 3848
rect 1607 3814 1623 3848
rect 1666 3846 1700 3862
rect 138 3750 172 3766
rect 215 3718 231 3752
rect 1607 3718 1623 3752
rect 1666 3704 1700 3720
rect 138 3608 172 3624
rect 215 3622 231 3656
rect 1607 3622 1623 3656
rect 1666 3654 1700 3670
rect 138 3558 172 3574
rect 215 3526 231 3560
rect 1607 3526 1623 3560
rect 1666 3512 1700 3528
rect 138 3416 172 3432
rect 215 3430 231 3464
rect 1607 3430 1623 3464
rect 1666 3462 1700 3478
rect 138 3366 172 3382
rect 215 3334 231 3368
rect 1607 3334 1623 3368
rect 1666 3320 1700 3336
rect 138 3224 172 3240
rect 215 3238 231 3272
rect 1607 3238 1623 3272
rect 1666 3270 1700 3286
rect 138 3174 172 3190
rect 215 3142 231 3176
rect 1607 3142 1623 3176
rect 1666 3128 1700 3144
rect 138 3032 172 3048
rect 215 3046 231 3080
rect 1607 3046 1623 3080
rect 1666 3078 1700 3094
rect 138 2982 172 2998
rect 215 2950 231 2984
rect 1607 2950 1623 2984
rect 1666 2936 1700 2952
rect 138 2840 172 2856
rect 215 2854 231 2888
rect 1607 2854 1623 2888
rect 1666 2886 1700 2902
rect 138 2790 172 2806
rect 215 2758 231 2792
rect 1607 2758 1623 2792
rect 1666 2744 1700 2760
rect 138 2648 172 2664
rect 215 2662 231 2696
rect 1607 2662 1623 2696
rect 1666 2694 1700 2710
rect 138 2598 172 2614
rect 215 2566 231 2600
rect 1607 2566 1623 2600
rect 1666 2552 1700 2568
rect 138 2456 172 2472
rect 215 2470 231 2504
rect 1607 2470 1623 2504
rect 1666 2502 1700 2518
rect 138 2406 172 2422
rect 215 2374 231 2408
rect 1607 2374 1623 2408
rect 1666 2360 1700 2376
rect 138 2264 172 2280
rect 215 2278 231 2312
rect 1607 2278 1623 2312
rect 1666 2310 1700 2326
rect 138 2214 172 2230
rect 215 2182 231 2216
rect 1607 2182 1623 2216
rect 1666 2168 1700 2184
rect 138 2072 172 2088
rect 215 2086 231 2120
rect 1607 2086 1623 2120
rect 1666 2118 1700 2134
rect 138 2022 172 2038
rect 215 1990 231 2024
rect 1607 1990 1623 2024
rect 1666 1976 1700 1992
rect 138 1880 172 1896
rect 215 1894 231 1928
rect 1607 1894 1623 1928
rect 1666 1926 1700 1942
rect 138 1830 172 1846
rect 215 1798 231 1832
rect 1607 1798 1623 1832
rect 1666 1784 1700 1800
rect 138 1688 172 1704
rect 215 1702 231 1736
rect 1607 1702 1623 1736
rect 1666 1734 1700 1750
rect 138 1638 172 1654
rect 215 1606 231 1640
rect 1607 1606 1623 1640
rect 1666 1592 1700 1608
rect 138 1496 172 1512
rect 215 1510 231 1544
rect 1607 1510 1623 1544
rect 1666 1542 1700 1558
rect 138 1446 172 1462
rect 215 1414 231 1448
rect 1607 1414 1623 1448
rect 1666 1400 1700 1416
rect 138 1304 172 1320
rect 215 1318 231 1352
rect 1607 1318 1623 1352
rect 1666 1350 1700 1366
rect 138 1254 172 1270
rect 215 1222 231 1256
rect 1607 1222 1623 1256
rect 1666 1208 1700 1224
rect 138 1112 172 1128
rect 215 1126 231 1160
rect 1607 1126 1623 1160
rect 1666 1158 1700 1174
rect 138 1062 172 1078
rect 215 1030 231 1064
rect 1607 1030 1623 1064
rect 1666 1016 1700 1032
rect 138 920 172 936
rect 215 934 231 968
rect 1607 934 1623 968
rect 1666 966 1700 982
rect 138 870 172 886
rect 215 838 231 872
rect 1607 838 1623 872
rect 1666 824 1700 840
rect 138 728 172 744
rect 215 742 231 776
rect 1607 742 1623 776
rect 1666 774 1700 790
rect 138 678 172 694
rect 215 646 231 680
rect 1607 646 1623 680
rect 1666 632 1700 648
rect 215 550 231 584
rect 1607 550 1623 584
rect 1666 582 1700 598
rect 36 470 70 532
rect 1768 470 1802 532
rect 36 436 132 470
rect 1706 436 1802 470
<< viali >>
rect 231 44168 1607 44202
rect 138 44120 172 44154
rect 231 44072 1607 44106
rect 1666 44024 1700 44058
rect 231 43976 1607 44010
rect 138 43928 172 43962
rect 231 43880 1607 43914
rect 1666 43832 1700 43866
rect 231 43784 1607 43818
rect 138 43736 172 43770
rect 231 43688 1607 43722
rect 1666 43640 1700 43674
rect 231 43592 1607 43626
rect 138 43544 172 43578
rect 231 43496 1607 43530
rect 1666 43448 1700 43482
rect 231 43400 1607 43434
rect 138 43352 172 43386
rect 231 43304 1607 43338
rect 1666 43256 1700 43290
rect 231 43208 1607 43242
rect 138 43160 172 43194
rect 231 43112 1607 43146
rect 1666 43064 1700 43098
rect 231 43016 1607 43050
rect 138 42968 172 43002
rect 231 42920 1607 42954
rect 1666 42872 1700 42906
rect 231 42824 1607 42858
rect 138 42776 172 42810
rect 231 42728 1607 42762
rect 1666 42680 1700 42714
rect 231 42632 1607 42666
rect 138 42584 172 42618
rect 231 42536 1607 42570
rect 1666 42488 1700 42522
rect 231 42440 1607 42474
rect 138 42392 172 42426
rect 231 42344 1607 42378
rect 1666 42296 1700 42330
rect 231 42248 1607 42282
rect 138 42200 172 42234
rect 231 42152 1607 42186
rect 1666 42104 1700 42138
rect 231 42056 1607 42090
rect 138 42008 172 42042
rect 231 41960 1607 41994
rect 1666 41912 1700 41946
rect 231 41864 1607 41898
rect 138 41816 172 41850
rect 231 41768 1607 41802
rect 1666 41720 1700 41754
rect 231 41672 1607 41706
rect 138 41624 172 41658
rect 231 41576 1607 41610
rect 1666 41528 1700 41562
rect 231 41480 1607 41514
rect 138 41432 172 41466
rect 231 41384 1607 41418
rect 1666 41336 1700 41370
rect 231 41288 1607 41322
rect 138 41240 172 41274
rect 231 41192 1607 41226
rect 1666 41144 1700 41178
rect 231 41096 1607 41130
rect 138 41048 172 41082
rect 231 41000 1607 41034
rect 1666 40952 1700 40986
rect 231 40904 1607 40938
rect 138 40856 172 40890
rect 231 40808 1607 40842
rect 1666 40760 1700 40794
rect 231 40712 1607 40746
rect 138 40664 172 40698
rect 231 40616 1607 40650
rect 1666 40568 1700 40602
rect 231 40520 1607 40554
rect 138 40472 172 40506
rect 231 40424 1607 40458
rect 1666 40376 1700 40410
rect 231 40328 1607 40362
rect 138 40280 172 40314
rect 231 40232 1607 40266
rect 1666 40184 1700 40218
rect 231 40136 1607 40170
rect 138 40088 172 40122
rect 231 40040 1607 40074
rect 1666 39992 1700 40026
rect 231 39944 1607 39978
rect 138 39896 172 39930
rect 231 39848 1607 39882
rect 1666 39800 1700 39834
rect 231 39752 1607 39786
rect 138 39704 172 39738
rect 231 39656 1607 39690
rect 1666 39608 1700 39642
rect 231 39560 1607 39594
rect 138 39512 172 39546
rect 231 39464 1607 39498
rect 1666 39416 1700 39450
rect 231 39368 1607 39402
rect 138 39320 172 39354
rect 231 39272 1607 39306
rect 1666 39224 1700 39258
rect 231 39176 1607 39210
rect 138 39128 172 39162
rect 231 39080 1607 39114
rect 1666 39032 1700 39066
rect 231 38984 1607 39018
rect 138 38936 172 38970
rect 231 38888 1607 38922
rect 1666 38840 1700 38874
rect 231 38792 1607 38826
rect 138 38744 172 38778
rect 231 38696 1607 38730
rect 1666 38648 1700 38682
rect 231 38600 1607 38634
rect 138 38552 172 38586
rect 231 38504 1607 38538
rect 1666 38456 1700 38490
rect 231 38408 1607 38442
rect 138 38360 172 38394
rect 231 38312 1607 38346
rect 1666 38264 1700 38298
rect 231 38216 1607 38250
rect 138 38168 172 38202
rect 231 38120 1607 38154
rect 1666 38072 1700 38106
rect 231 38024 1607 38058
rect 138 37976 172 38010
rect 231 37928 1607 37962
rect 1666 37880 1700 37914
rect 231 37832 1607 37866
rect 138 37784 172 37818
rect 231 37736 1607 37770
rect 1666 37688 1700 37722
rect 231 37640 1607 37674
rect 138 37592 172 37626
rect 231 37544 1607 37578
rect 1666 37496 1700 37530
rect 231 37448 1607 37482
rect 138 37400 172 37434
rect 231 37352 1607 37386
rect 1666 37304 1700 37338
rect 231 37256 1607 37290
rect 138 37208 172 37242
rect 231 37160 1607 37194
rect 1666 37112 1700 37146
rect 231 37064 1607 37098
rect 138 37016 172 37050
rect 231 36968 1607 37002
rect 1666 36920 1700 36954
rect 231 36872 1607 36906
rect 138 36824 172 36858
rect 231 36776 1607 36810
rect 1666 36728 1700 36762
rect 231 36680 1607 36714
rect 138 36632 172 36666
rect 231 36584 1607 36618
rect 1666 36536 1700 36570
rect 231 36488 1607 36522
rect 138 36440 172 36474
rect 231 36392 1607 36426
rect 1666 36344 1700 36378
rect 231 36296 1607 36330
rect 138 36248 172 36282
rect 231 36200 1607 36234
rect 1666 36152 1700 36186
rect 231 36104 1607 36138
rect 138 36056 172 36090
rect 231 36008 1607 36042
rect 1666 35960 1700 35994
rect 231 35912 1607 35946
rect 138 35864 172 35898
rect 231 35816 1607 35850
rect 1666 35768 1700 35802
rect 231 35720 1607 35754
rect 138 35672 172 35706
rect 231 35624 1607 35658
rect 1666 35576 1700 35610
rect 231 35528 1607 35562
rect 138 35480 172 35514
rect 231 35432 1607 35466
rect 1666 35384 1700 35418
rect 231 35336 1607 35370
rect 138 35288 172 35322
rect 231 35240 1607 35274
rect 1666 35192 1700 35226
rect 231 35144 1607 35178
rect 138 35096 172 35130
rect 231 35048 1607 35082
rect 1666 35000 1700 35034
rect 231 34952 1607 34986
rect 138 34904 172 34938
rect 231 34856 1607 34890
rect 1666 34808 1700 34842
rect 231 34760 1607 34794
rect 138 34712 172 34746
rect 231 34664 1607 34698
rect 1666 34616 1700 34650
rect 231 34568 1607 34602
rect 138 34520 172 34554
rect 231 34472 1607 34506
rect 1666 34424 1700 34458
rect 231 34376 1607 34410
rect 138 34328 172 34362
rect 231 34280 1607 34314
rect 1666 34232 1700 34266
rect 231 34184 1607 34218
rect 138 34136 172 34170
rect 231 34088 1607 34122
rect 1666 34040 1700 34074
rect 231 33992 1607 34026
rect 138 33944 172 33978
rect 231 33896 1607 33930
rect 1666 33848 1700 33882
rect 231 33800 1607 33834
rect 138 33752 172 33786
rect 231 33704 1607 33738
rect 1666 33656 1700 33690
rect 231 33608 1607 33642
rect 138 33560 172 33594
rect 231 33512 1607 33546
rect 1666 33464 1700 33498
rect 231 33416 1607 33450
rect 138 33368 172 33402
rect 231 33320 1607 33354
rect 1666 33272 1700 33306
rect 231 33224 1607 33258
rect 138 33176 172 33210
rect 231 33128 1607 33162
rect 1666 33080 1700 33114
rect 231 33032 1607 33066
rect 138 32984 172 33018
rect 231 32936 1607 32970
rect 1666 32888 1700 32922
rect 231 32840 1607 32874
rect 138 32792 172 32826
rect 231 32744 1607 32778
rect 1666 32696 1700 32730
rect 231 32648 1607 32682
rect 138 32600 172 32634
rect 231 32552 1607 32586
rect 1666 32504 1700 32538
rect 231 32456 1607 32490
rect 138 32408 172 32442
rect 231 32360 1607 32394
rect 1666 32312 1700 32346
rect 231 32264 1607 32298
rect 138 32216 172 32250
rect 231 32168 1607 32202
rect 1666 32120 1700 32154
rect 231 32072 1607 32106
rect 138 32024 172 32058
rect 231 31976 1607 32010
rect 1666 31928 1700 31962
rect 231 31880 1607 31914
rect 138 31832 172 31866
rect 231 31784 1607 31818
rect 1666 31736 1700 31770
rect 231 31688 1607 31722
rect 138 31640 172 31674
rect 231 31592 1607 31626
rect 1666 31544 1700 31578
rect 231 31496 1607 31530
rect 138 31448 172 31482
rect 231 31400 1607 31434
rect 1666 31352 1700 31386
rect 231 31304 1607 31338
rect 138 31256 172 31290
rect 231 31208 1607 31242
rect 1666 31160 1700 31194
rect 231 31112 1607 31146
rect 138 31064 172 31098
rect 231 31016 1607 31050
rect 1666 30968 1700 31002
rect 231 30920 1607 30954
rect 138 30872 172 30906
rect 231 30824 1607 30858
rect 1666 30776 1700 30810
rect 231 30728 1607 30762
rect 138 30680 172 30714
rect 231 30632 1607 30666
rect 1666 30584 1700 30618
rect 231 30536 1607 30570
rect 138 30488 172 30522
rect 231 30440 1607 30474
rect 1666 30392 1700 30426
rect 231 30344 1607 30378
rect 138 30296 172 30330
rect 231 30248 1607 30282
rect 1666 30200 1700 30234
rect 231 30152 1607 30186
rect 138 30104 172 30138
rect 231 30056 1607 30090
rect 1666 30008 1700 30042
rect 231 29960 1607 29994
rect 138 29912 172 29946
rect 231 29864 1607 29898
rect 1666 29816 1700 29850
rect 231 29768 1607 29802
rect 138 29720 172 29754
rect 231 29672 1607 29706
rect 1666 29624 1700 29658
rect 231 29576 1607 29610
rect 138 29528 172 29562
rect 231 29480 1607 29514
rect 1666 29432 1700 29466
rect 231 29384 1607 29418
rect 138 29336 172 29370
rect 231 29288 1607 29322
rect 1666 29240 1700 29274
rect 231 29192 1607 29226
rect 138 29144 172 29178
rect 231 29096 1607 29130
rect 1666 29048 1700 29082
rect 231 29000 1607 29034
rect 138 28952 172 28986
rect 231 28904 1607 28938
rect 1666 28856 1700 28890
rect 231 28808 1607 28842
rect 138 28760 172 28794
rect 231 28712 1607 28746
rect 1666 28664 1700 28698
rect 231 28616 1607 28650
rect 138 28568 172 28602
rect 231 28520 1607 28554
rect 1666 28472 1700 28506
rect 231 28424 1607 28458
rect 138 28376 172 28410
rect 231 28328 1607 28362
rect 1666 28280 1700 28314
rect 231 28232 1607 28266
rect 138 28184 172 28218
rect 231 28136 1607 28170
rect 1666 28088 1700 28122
rect 231 28040 1607 28074
rect 138 27992 172 28026
rect 231 27944 1607 27978
rect 1666 27896 1700 27930
rect 231 27848 1607 27882
rect 138 27800 172 27834
rect 231 27752 1607 27786
rect 1666 27704 1700 27738
rect 231 27656 1607 27690
rect 138 27608 172 27642
rect 231 27560 1607 27594
rect 1666 27512 1700 27546
rect 231 27464 1607 27498
rect 138 27416 172 27450
rect 231 27368 1607 27402
rect 1666 27320 1700 27354
rect 231 27272 1607 27306
rect 138 27224 172 27258
rect 231 27176 1607 27210
rect 1666 27128 1700 27162
rect 231 27080 1607 27114
rect 138 27032 172 27066
rect 231 26984 1607 27018
rect 1666 26936 1700 26970
rect 231 26888 1607 26922
rect 138 26840 172 26874
rect 231 26792 1607 26826
rect 1666 26744 1700 26778
rect 231 26696 1607 26730
rect 138 26648 172 26682
rect 231 26600 1607 26634
rect 1666 26552 1700 26586
rect 231 26504 1607 26538
rect 138 26456 172 26490
rect 231 26408 1607 26442
rect 1666 26360 1700 26394
rect 231 26312 1607 26346
rect 138 26264 172 26298
rect 231 26216 1607 26250
rect 1666 26168 1700 26202
rect 231 26120 1607 26154
rect 138 26072 172 26106
rect 231 26024 1607 26058
rect 1666 25976 1700 26010
rect 231 25928 1607 25962
rect 138 25880 172 25914
rect 231 25832 1607 25866
rect 1666 25784 1700 25818
rect 231 25736 1607 25770
rect 138 25688 172 25722
rect 231 25640 1607 25674
rect 1666 25592 1700 25626
rect 231 25544 1607 25578
rect 138 25496 172 25530
rect 231 25448 1607 25482
rect 1666 25400 1700 25434
rect 231 25352 1607 25386
rect 138 25304 172 25338
rect 231 25256 1607 25290
rect 1666 25208 1700 25242
rect 231 25160 1607 25194
rect 138 25112 172 25146
rect 231 25064 1607 25098
rect 1666 25016 1700 25050
rect 231 24968 1607 25002
rect 138 24920 172 24954
rect 231 24872 1607 24906
rect 1666 24824 1700 24858
rect 231 24776 1607 24810
rect 138 24728 172 24762
rect 231 24680 1607 24714
rect 1666 24632 1700 24666
rect 231 24584 1607 24618
rect 138 24536 172 24570
rect 231 24488 1607 24522
rect 1666 24440 1700 24474
rect 231 24392 1607 24426
rect 138 24344 172 24378
rect 231 24296 1607 24330
rect 1666 24248 1700 24282
rect 231 24200 1607 24234
rect 138 24152 172 24186
rect 231 24104 1607 24138
rect 1666 24056 1700 24090
rect 231 24008 1607 24042
rect 138 23960 172 23994
rect 231 23912 1607 23946
rect 1666 23864 1700 23898
rect 231 23816 1607 23850
rect 138 23768 172 23802
rect 231 23720 1607 23754
rect 1666 23672 1700 23706
rect 231 23624 1607 23658
rect 138 23576 172 23610
rect 231 23528 1607 23562
rect 1666 23480 1700 23514
rect 231 23432 1607 23466
rect 138 23384 172 23418
rect 231 23336 1607 23370
rect 1666 23288 1700 23322
rect 231 23240 1607 23274
rect 138 23192 172 23226
rect 231 23144 1607 23178
rect 1666 23096 1700 23130
rect 231 23048 1607 23082
rect 340 21986 870 22768
rect 231 21670 1607 21704
rect 138 21622 172 21656
rect 231 21574 1607 21608
rect 1666 21526 1700 21560
rect 231 21478 1607 21512
rect 138 21430 172 21464
rect 231 21382 1607 21416
rect 1666 21334 1700 21368
rect 231 21286 1607 21320
rect 138 21238 172 21272
rect 231 21190 1607 21224
rect 1666 21142 1700 21176
rect 231 21094 1607 21128
rect 138 21046 172 21080
rect 231 20998 1607 21032
rect 1666 20950 1700 20984
rect 231 20902 1607 20936
rect 138 20854 172 20888
rect 231 20806 1607 20840
rect 1666 20758 1700 20792
rect 231 20710 1607 20744
rect 138 20662 172 20696
rect 231 20614 1607 20648
rect 1666 20566 1700 20600
rect 231 20518 1607 20552
rect 138 20470 172 20504
rect 231 20422 1607 20456
rect 1666 20374 1700 20408
rect 231 20326 1607 20360
rect 138 20278 172 20312
rect 231 20230 1607 20264
rect 1666 20182 1700 20216
rect 231 20134 1607 20168
rect 138 20086 172 20120
rect 231 20038 1607 20072
rect 1666 19990 1700 20024
rect 231 19942 1607 19976
rect 138 19894 172 19928
rect 231 19846 1607 19880
rect 1666 19798 1700 19832
rect 231 19750 1607 19784
rect 138 19702 172 19736
rect 231 19654 1607 19688
rect 1666 19606 1700 19640
rect 231 19558 1607 19592
rect 138 19510 172 19544
rect 231 19462 1607 19496
rect 1666 19414 1700 19448
rect 231 19366 1607 19400
rect 138 19318 172 19352
rect 231 19270 1607 19304
rect 1666 19222 1700 19256
rect 231 19174 1607 19208
rect 138 19126 172 19160
rect 231 19078 1607 19112
rect 1666 19030 1700 19064
rect 231 18982 1607 19016
rect 138 18934 172 18968
rect 231 18886 1607 18920
rect 1666 18838 1700 18872
rect 231 18790 1607 18824
rect 138 18742 172 18776
rect 231 18694 1607 18728
rect 1666 18646 1700 18680
rect 231 18598 1607 18632
rect 138 18550 172 18584
rect 231 18502 1607 18536
rect 1666 18454 1700 18488
rect 231 18406 1607 18440
rect 138 18358 172 18392
rect 231 18310 1607 18344
rect 1666 18262 1700 18296
rect 231 18214 1607 18248
rect 138 18166 172 18200
rect 231 18118 1607 18152
rect 1666 18070 1700 18104
rect 231 18022 1607 18056
rect 138 17974 172 18008
rect 231 17926 1607 17960
rect 1666 17878 1700 17912
rect 231 17830 1607 17864
rect 138 17782 172 17816
rect 231 17734 1607 17768
rect 1666 17686 1700 17720
rect 231 17638 1607 17672
rect 138 17590 172 17624
rect 231 17542 1607 17576
rect 1666 17494 1700 17528
rect 231 17446 1607 17480
rect 138 17398 172 17432
rect 231 17350 1607 17384
rect 1666 17302 1700 17336
rect 231 17254 1607 17288
rect 138 17206 172 17240
rect 231 17158 1607 17192
rect 1666 17110 1700 17144
rect 231 17062 1607 17096
rect 138 17014 172 17048
rect 231 16966 1607 17000
rect 1666 16918 1700 16952
rect 231 16870 1607 16904
rect 138 16822 172 16856
rect 231 16774 1607 16808
rect 1666 16726 1700 16760
rect 231 16678 1607 16712
rect 138 16630 172 16664
rect 231 16582 1607 16616
rect 1666 16534 1700 16568
rect 231 16486 1607 16520
rect 138 16438 172 16472
rect 231 16390 1607 16424
rect 1666 16342 1700 16376
rect 231 16294 1607 16328
rect 138 16246 172 16280
rect 231 16198 1607 16232
rect 1666 16150 1700 16184
rect 231 16102 1607 16136
rect 138 16054 172 16088
rect 231 16006 1607 16040
rect 1666 15958 1700 15992
rect 231 15910 1607 15944
rect 138 15862 172 15896
rect 231 15814 1607 15848
rect 1666 15766 1700 15800
rect 231 15718 1607 15752
rect 138 15670 172 15704
rect 231 15622 1607 15656
rect 1666 15574 1700 15608
rect 231 15526 1607 15560
rect 138 15478 172 15512
rect 231 15430 1607 15464
rect 1666 15382 1700 15416
rect 231 15334 1607 15368
rect 138 15286 172 15320
rect 231 15238 1607 15272
rect 1666 15190 1700 15224
rect 231 15142 1607 15176
rect 138 15094 172 15128
rect 231 15046 1607 15080
rect 1666 14998 1700 15032
rect 231 14950 1607 14984
rect 138 14902 172 14936
rect 231 14854 1607 14888
rect 1666 14806 1700 14840
rect 231 14758 1607 14792
rect 138 14710 172 14744
rect 231 14662 1607 14696
rect 1666 14614 1700 14648
rect 231 14566 1607 14600
rect 138 14518 172 14552
rect 231 14470 1607 14504
rect 1666 14422 1700 14456
rect 231 14374 1607 14408
rect 138 14326 172 14360
rect 231 14278 1607 14312
rect 1666 14230 1700 14264
rect 231 14182 1607 14216
rect 138 14134 172 14168
rect 231 14086 1607 14120
rect 1666 14038 1700 14072
rect 231 13990 1607 14024
rect 138 13942 172 13976
rect 231 13894 1607 13928
rect 1666 13846 1700 13880
rect 231 13798 1607 13832
rect 138 13750 172 13784
rect 231 13702 1607 13736
rect 1666 13654 1700 13688
rect 231 13606 1607 13640
rect 138 13558 172 13592
rect 231 13510 1607 13544
rect 1666 13462 1700 13496
rect 231 13414 1607 13448
rect 138 13366 172 13400
rect 231 13318 1607 13352
rect 1666 13270 1700 13304
rect 231 13222 1607 13256
rect 138 13174 172 13208
rect 231 13126 1607 13160
rect 1666 13078 1700 13112
rect 231 13030 1607 13064
rect 138 12982 172 13016
rect 231 12934 1607 12968
rect 1666 12886 1700 12920
rect 231 12838 1607 12872
rect 138 12790 172 12824
rect 231 12742 1607 12776
rect 1666 12694 1700 12728
rect 231 12646 1607 12680
rect 138 12598 172 12632
rect 231 12550 1607 12584
rect 1666 12502 1700 12536
rect 231 12454 1607 12488
rect 138 12406 172 12440
rect 231 12358 1607 12392
rect 1666 12310 1700 12344
rect 231 12262 1607 12296
rect 138 12214 172 12248
rect 231 12166 1607 12200
rect 1666 12118 1700 12152
rect 231 12070 1607 12104
rect 138 12022 172 12056
rect 231 11974 1607 12008
rect 1666 11926 1700 11960
rect 231 11878 1607 11912
rect 138 11830 172 11864
rect 231 11782 1607 11816
rect 1666 11734 1700 11768
rect 231 11686 1607 11720
rect 138 11638 172 11672
rect 231 11590 1607 11624
rect 1666 11542 1700 11576
rect 231 11494 1607 11528
rect 138 11446 172 11480
rect 231 11398 1607 11432
rect 1666 11350 1700 11384
rect 231 11302 1607 11336
rect 138 11254 172 11288
rect 231 11206 1607 11240
rect 1666 11158 1700 11192
rect 231 11110 1607 11144
rect 138 11062 172 11096
rect 231 11014 1607 11048
rect 1666 10966 1700 11000
rect 231 10918 1607 10952
rect 138 10870 172 10904
rect 231 10822 1607 10856
rect 1666 10774 1700 10808
rect 231 10726 1607 10760
rect 138 10678 172 10712
rect 231 10630 1607 10664
rect 1666 10582 1700 10616
rect 231 10534 1607 10568
rect 138 10486 172 10520
rect 231 10438 1607 10472
rect 1666 10390 1700 10424
rect 231 10342 1607 10376
rect 138 10294 172 10328
rect 231 10246 1607 10280
rect 1666 10198 1700 10232
rect 231 10150 1607 10184
rect 138 10102 172 10136
rect 231 10054 1607 10088
rect 1666 10006 1700 10040
rect 231 9958 1607 9992
rect 138 9910 172 9944
rect 231 9862 1607 9896
rect 1666 9814 1700 9848
rect 231 9766 1607 9800
rect 138 9718 172 9752
rect 231 9670 1607 9704
rect 1666 9622 1700 9656
rect 231 9574 1607 9608
rect 138 9526 172 9560
rect 231 9478 1607 9512
rect 1666 9430 1700 9464
rect 231 9382 1607 9416
rect 138 9334 172 9368
rect 231 9286 1607 9320
rect 1666 9238 1700 9272
rect 231 9190 1607 9224
rect 138 9142 172 9176
rect 231 9094 1607 9128
rect 1666 9046 1700 9080
rect 231 8998 1607 9032
rect 138 8950 172 8984
rect 231 8902 1607 8936
rect 1666 8854 1700 8888
rect 231 8806 1607 8840
rect 138 8758 172 8792
rect 231 8710 1607 8744
rect 1666 8662 1700 8696
rect 231 8614 1607 8648
rect 138 8566 172 8600
rect 231 8518 1607 8552
rect 1666 8470 1700 8504
rect 231 8422 1607 8456
rect 138 8374 172 8408
rect 231 8326 1607 8360
rect 1666 8278 1700 8312
rect 231 8230 1607 8264
rect 138 8182 172 8216
rect 231 8134 1607 8168
rect 1666 8086 1700 8120
rect 231 8038 1607 8072
rect 138 7990 172 8024
rect 231 7942 1607 7976
rect 1666 7894 1700 7928
rect 231 7846 1607 7880
rect 138 7798 172 7832
rect 231 7750 1607 7784
rect 1666 7702 1700 7736
rect 231 7654 1607 7688
rect 138 7606 172 7640
rect 231 7558 1607 7592
rect 1666 7510 1700 7544
rect 231 7462 1607 7496
rect 138 7414 172 7448
rect 231 7366 1607 7400
rect 1666 7318 1700 7352
rect 231 7270 1607 7304
rect 138 7222 172 7256
rect 231 7174 1607 7208
rect 1666 7126 1700 7160
rect 231 7078 1607 7112
rect 138 7030 172 7064
rect 231 6982 1607 7016
rect 1666 6934 1700 6968
rect 231 6886 1607 6920
rect 138 6838 172 6872
rect 231 6790 1607 6824
rect 1666 6742 1700 6776
rect 231 6694 1607 6728
rect 138 6646 172 6680
rect 231 6598 1607 6632
rect 1666 6550 1700 6584
rect 231 6502 1607 6536
rect 138 6454 172 6488
rect 231 6406 1607 6440
rect 1666 6358 1700 6392
rect 231 6310 1607 6344
rect 138 6262 172 6296
rect 231 6214 1607 6248
rect 1666 6166 1700 6200
rect 231 6118 1607 6152
rect 138 6070 172 6104
rect 231 6022 1607 6056
rect 1666 5974 1700 6008
rect 231 5926 1607 5960
rect 138 5878 172 5912
rect 231 5830 1607 5864
rect 1666 5782 1700 5816
rect 231 5734 1607 5768
rect 138 5686 172 5720
rect 231 5638 1607 5672
rect 1666 5590 1700 5624
rect 231 5542 1607 5576
rect 138 5494 172 5528
rect 231 5446 1607 5480
rect 1666 5398 1700 5432
rect 231 5350 1607 5384
rect 138 5302 172 5336
rect 231 5254 1607 5288
rect 1666 5206 1700 5240
rect 231 5158 1607 5192
rect 138 5110 172 5144
rect 231 5062 1607 5096
rect 1666 5014 1700 5048
rect 231 4966 1607 5000
rect 138 4918 172 4952
rect 231 4870 1607 4904
rect 1666 4822 1700 4856
rect 231 4774 1607 4808
rect 138 4726 172 4760
rect 231 4678 1607 4712
rect 1666 4630 1700 4664
rect 231 4582 1607 4616
rect 138 4534 172 4568
rect 231 4486 1607 4520
rect 1666 4438 1700 4472
rect 231 4390 1607 4424
rect 138 4342 172 4376
rect 231 4294 1607 4328
rect 1666 4246 1700 4280
rect 231 4198 1607 4232
rect 138 4150 172 4184
rect 231 4102 1607 4136
rect 1666 4054 1700 4088
rect 231 4006 1607 4040
rect 138 3958 172 3992
rect 231 3910 1607 3944
rect 1666 3862 1700 3896
rect 231 3814 1607 3848
rect 138 3766 172 3800
rect 231 3718 1607 3752
rect 1666 3670 1700 3704
rect 231 3622 1607 3656
rect 138 3574 172 3608
rect 231 3526 1607 3560
rect 1666 3478 1700 3512
rect 231 3430 1607 3464
rect 138 3382 172 3416
rect 231 3334 1607 3368
rect 1666 3286 1700 3320
rect 231 3238 1607 3272
rect 138 3190 172 3224
rect 231 3142 1607 3176
rect 1666 3094 1700 3128
rect 231 3046 1607 3080
rect 138 2998 172 3032
rect 231 2950 1607 2984
rect 1666 2902 1700 2936
rect 231 2854 1607 2888
rect 138 2806 172 2840
rect 231 2758 1607 2792
rect 1666 2710 1700 2744
rect 231 2662 1607 2696
rect 138 2614 172 2648
rect 231 2566 1607 2600
rect 1666 2518 1700 2552
rect 231 2470 1607 2504
rect 138 2422 172 2456
rect 231 2374 1607 2408
rect 1666 2326 1700 2360
rect 231 2278 1607 2312
rect 138 2230 172 2264
rect 231 2182 1607 2216
rect 1666 2134 1700 2168
rect 231 2086 1607 2120
rect 138 2038 172 2072
rect 231 1990 1607 2024
rect 1666 1942 1700 1976
rect 231 1894 1607 1928
rect 138 1846 172 1880
rect 231 1798 1607 1832
rect 1666 1750 1700 1784
rect 231 1702 1607 1736
rect 138 1654 172 1688
rect 231 1606 1607 1640
rect 1666 1558 1700 1592
rect 231 1510 1607 1544
rect 138 1462 172 1496
rect 231 1414 1607 1448
rect 1666 1366 1700 1400
rect 231 1318 1607 1352
rect 138 1270 172 1304
rect 231 1222 1607 1256
rect 1666 1174 1700 1208
rect 231 1126 1607 1160
rect 138 1078 172 1112
rect 231 1030 1607 1064
rect 1666 982 1700 1016
rect 231 934 1607 968
rect 138 886 172 920
rect 231 838 1607 872
rect 1666 790 1700 824
rect 231 742 1607 776
rect 138 694 172 728
rect 231 646 1607 680
rect 1666 598 1700 632
rect 231 550 1607 584
<< metal1 >>
rect 122 45072 132 45126
rect 1706 45072 1716 45126
rect 132 44154 178 45072
rect 342 44208 352 44218
rect 219 44202 352 44208
rect 858 44208 868 44218
rect 858 44202 1619 44208
rect 219 44168 231 44202
rect 1607 44168 1619 44202
rect 219 44162 352 44168
rect 132 44120 138 44154
rect 172 44120 178 44154
rect 342 44152 352 44162
rect 858 44162 1619 44168
rect 858 44152 868 44162
rect 132 43962 178 44120
rect 970 44112 980 44122
rect 219 44106 980 44112
rect 1490 44112 1500 44122
rect 1490 44106 1619 44112
rect 219 44072 231 44106
rect 1607 44072 1619 44106
rect 219 44066 980 44072
rect 970 44056 980 44066
rect 1490 44066 1619 44072
rect 1490 44056 1500 44066
rect 1660 44058 1706 45072
rect 342 44016 352 44026
rect 219 44010 352 44016
rect 858 44016 868 44026
rect 1660 44024 1666 44058
rect 1700 44024 1706 44058
rect 858 44010 1619 44016
rect 219 43976 231 44010
rect 1607 43976 1619 44010
rect 219 43970 352 43976
rect 132 43928 138 43962
rect 172 43928 178 43962
rect 342 43960 352 43970
rect 858 43970 1619 43976
rect 858 43960 868 43970
rect 132 43770 178 43928
rect 970 43920 980 43930
rect 219 43914 980 43920
rect 1490 43920 1500 43930
rect 1490 43914 1619 43920
rect 219 43880 231 43914
rect 1607 43880 1619 43914
rect 219 43874 980 43880
rect 970 43864 980 43874
rect 1490 43874 1619 43880
rect 1490 43864 1500 43874
rect 1660 43866 1706 44024
rect 342 43824 352 43834
rect 219 43818 352 43824
rect 858 43824 868 43834
rect 1660 43832 1666 43866
rect 1700 43832 1706 43866
rect 858 43818 1619 43824
rect 219 43784 231 43818
rect 1607 43784 1619 43818
rect 219 43778 352 43784
rect 132 43736 138 43770
rect 172 43736 178 43770
rect 342 43768 352 43778
rect 858 43778 1619 43784
rect 858 43768 868 43778
rect 132 43578 178 43736
rect 970 43728 980 43738
rect 219 43722 980 43728
rect 1490 43728 1500 43738
rect 1490 43722 1619 43728
rect 219 43688 231 43722
rect 1607 43688 1619 43722
rect 219 43682 980 43688
rect 970 43672 980 43682
rect 1490 43682 1619 43688
rect 1490 43672 1500 43682
rect 1660 43674 1706 43832
rect 342 43632 352 43642
rect 219 43626 352 43632
rect 858 43632 868 43642
rect 1660 43640 1666 43674
rect 1700 43640 1706 43674
rect 858 43626 1619 43632
rect 219 43592 231 43626
rect 1607 43592 1619 43626
rect 219 43586 352 43592
rect 132 43544 138 43578
rect 172 43544 178 43578
rect 342 43576 352 43586
rect 858 43586 1619 43592
rect 858 43576 868 43586
rect 132 43386 178 43544
rect 970 43536 980 43546
rect 219 43530 980 43536
rect 1490 43536 1500 43546
rect 1490 43530 1619 43536
rect 219 43496 231 43530
rect 1607 43496 1619 43530
rect 219 43490 980 43496
rect 970 43480 980 43490
rect 1490 43490 1619 43496
rect 1490 43480 1500 43490
rect 1660 43482 1706 43640
rect 342 43440 352 43450
rect 219 43434 352 43440
rect 858 43440 868 43450
rect 1660 43448 1666 43482
rect 1700 43448 1706 43482
rect 858 43434 1619 43440
rect 219 43400 231 43434
rect 1607 43400 1619 43434
rect 219 43394 352 43400
rect 132 43352 138 43386
rect 172 43352 178 43386
rect 342 43384 352 43394
rect 858 43394 1619 43400
rect 858 43384 868 43394
rect 132 43194 178 43352
rect 970 43344 980 43354
rect 219 43338 980 43344
rect 1490 43344 1500 43354
rect 1490 43338 1619 43344
rect 219 43304 231 43338
rect 1607 43304 1619 43338
rect 219 43298 980 43304
rect 970 43288 980 43298
rect 1490 43298 1619 43304
rect 1490 43288 1500 43298
rect 1660 43290 1706 43448
rect 342 43248 352 43258
rect 219 43242 352 43248
rect 858 43248 868 43258
rect 1660 43256 1666 43290
rect 1700 43256 1706 43290
rect 858 43242 1619 43248
rect 219 43208 231 43242
rect 1607 43208 1619 43242
rect 219 43202 352 43208
rect 132 43160 138 43194
rect 172 43160 178 43194
rect 342 43192 352 43202
rect 858 43202 1619 43208
rect 858 43192 868 43202
rect 132 43002 178 43160
rect 970 43152 980 43162
rect 219 43146 980 43152
rect 1490 43152 1500 43162
rect 1490 43146 1619 43152
rect 219 43112 231 43146
rect 1607 43112 1619 43146
rect 219 43106 980 43112
rect 970 43096 980 43106
rect 1490 43106 1619 43112
rect 1490 43096 1500 43106
rect 1660 43098 1706 43256
rect 342 43056 352 43066
rect 219 43050 352 43056
rect 858 43056 868 43066
rect 1660 43064 1666 43098
rect 1700 43064 1706 43098
rect 858 43050 1619 43056
rect 219 43016 231 43050
rect 1607 43016 1619 43050
rect 219 43010 352 43016
rect 132 42968 138 43002
rect 172 42968 178 43002
rect 342 43000 352 43010
rect 858 43010 1619 43016
rect 858 43000 868 43010
rect 132 42810 178 42968
rect 970 42960 980 42970
rect 219 42954 980 42960
rect 1490 42960 1500 42970
rect 1490 42954 1619 42960
rect 219 42920 231 42954
rect 1607 42920 1619 42954
rect 219 42914 980 42920
rect 970 42904 980 42914
rect 1490 42914 1619 42920
rect 1490 42904 1500 42914
rect 1660 42906 1706 43064
rect 342 42864 352 42874
rect 219 42858 352 42864
rect 858 42864 868 42874
rect 1660 42872 1666 42906
rect 1700 42872 1706 42906
rect 858 42858 1619 42864
rect 219 42824 231 42858
rect 1607 42824 1619 42858
rect 219 42818 352 42824
rect 132 42776 138 42810
rect 172 42776 178 42810
rect 342 42808 352 42818
rect 858 42818 1619 42824
rect 858 42808 868 42818
rect 132 42618 178 42776
rect 970 42768 980 42778
rect 219 42762 980 42768
rect 1490 42768 1500 42778
rect 1490 42762 1619 42768
rect 219 42728 231 42762
rect 1607 42728 1619 42762
rect 219 42722 980 42728
rect 970 42712 980 42722
rect 1490 42722 1619 42728
rect 1490 42712 1500 42722
rect 1660 42714 1706 42872
rect 342 42672 352 42682
rect 219 42666 352 42672
rect 858 42672 868 42682
rect 1660 42680 1666 42714
rect 1700 42680 1706 42714
rect 858 42666 1619 42672
rect 219 42632 231 42666
rect 1607 42632 1619 42666
rect 219 42626 352 42632
rect 132 42584 138 42618
rect 172 42584 178 42618
rect 342 42616 352 42626
rect 858 42626 1619 42632
rect 858 42616 868 42626
rect 132 42426 178 42584
rect 970 42576 980 42586
rect 219 42570 980 42576
rect 1490 42576 1500 42586
rect 1490 42570 1619 42576
rect 219 42536 231 42570
rect 1607 42536 1619 42570
rect 219 42530 980 42536
rect 970 42520 980 42530
rect 1490 42530 1619 42536
rect 1490 42520 1500 42530
rect 1660 42522 1706 42680
rect 342 42480 352 42490
rect 219 42474 352 42480
rect 858 42480 868 42490
rect 1660 42488 1666 42522
rect 1700 42488 1706 42522
rect 858 42474 1619 42480
rect 219 42440 231 42474
rect 1607 42440 1619 42474
rect 219 42434 352 42440
rect 132 42392 138 42426
rect 172 42392 178 42426
rect 342 42424 352 42434
rect 858 42434 1619 42440
rect 858 42424 868 42434
rect 132 42234 178 42392
rect 970 42384 980 42394
rect 219 42378 980 42384
rect 1490 42384 1500 42394
rect 1490 42378 1619 42384
rect 219 42344 231 42378
rect 1607 42344 1619 42378
rect 219 42338 980 42344
rect 970 42328 980 42338
rect 1490 42338 1619 42344
rect 1490 42328 1500 42338
rect 1660 42330 1706 42488
rect 342 42288 352 42298
rect 219 42282 352 42288
rect 858 42288 868 42298
rect 1660 42296 1666 42330
rect 1700 42296 1706 42330
rect 858 42282 1619 42288
rect 219 42248 231 42282
rect 1607 42248 1619 42282
rect 219 42242 352 42248
rect 132 42200 138 42234
rect 172 42200 178 42234
rect 342 42232 352 42242
rect 858 42242 1619 42248
rect 858 42232 868 42242
rect 132 42042 178 42200
rect 970 42192 980 42202
rect 219 42186 980 42192
rect 1490 42192 1500 42202
rect 1490 42186 1619 42192
rect 219 42152 231 42186
rect 1607 42152 1619 42186
rect 219 42146 980 42152
rect 970 42136 980 42146
rect 1490 42146 1619 42152
rect 1490 42136 1500 42146
rect 1660 42138 1706 42296
rect 342 42096 352 42106
rect 219 42090 352 42096
rect 858 42096 868 42106
rect 1660 42104 1666 42138
rect 1700 42104 1706 42138
rect 858 42090 1619 42096
rect 219 42056 231 42090
rect 1607 42056 1619 42090
rect 219 42050 352 42056
rect 132 42008 138 42042
rect 172 42008 178 42042
rect 342 42040 352 42050
rect 858 42050 1619 42056
rect 858 42040 868 42050
rect 132 41850 178 42008
rect 970 42000 980 42010
rect 219 41994 980 42000
rect 1490 42000 1500 42010
rect 1490 41994 1619 42000
rect 219 41960 231 41994
rect 1607 41960 1619 41994
rect 219 41954 980 41960
rect 970 41944 980 41954
rect 1490 41954 1619 41960
rect 1490 41944 1500 41954
rect 1660 41946 1706 42104
rect 342 41904 352 41914
rect 219 41898 352 41904
rect 858 41904 868 41914
rect 1660 41912 1666 41946
rect 1700 41912 1706 41946
rect 858 41898 1619 41904
rect 219 41864 231 41898
rect 1607 41864 1619 41898
rect 219 41858 352 41864
rect 132 41816 138 41850
rect 172 41816 178 41850
rect 342 41848 352 41858
rect 858 41858 1619 41864
rect 858 41848 868 41858
rect 132 41658 178 41816
rect 970 41808 980 41818
rect 219 41802 980 41808
rect 1490 41808 1500 41818
rect 1490 41802 1619 41808
rect 219 41768 231 41802
rect 1607 41768 1619 41802
rect 219 41762 980 41768
rect 970 41752 980 41762
rect 1490 41762 1619 41768
rect 1490 41752 1500 41762
rect 1660 41754 1706 41912
rect 342 41712 352 41722
rect 219 41706 352 41712
rect 858 41712 868 41722
rect 1660 41720 1666 41754
rect 1700 41720 1706 41754
rect 858 41706 1619 41712
rect 219 41672 231 41706
rect 1607 41672 1619 41706
rect 219 41666 352 41672
rect 132 41624 138 41658
rect 172 41624 178 41658
rect 342 41656 352 41666
rect 858 41666 1619 41672
rect 858 41656 868 41666
rect 132 41466 178 41624
rect 970 41616 980 41626
rect 219 41610 980 41616
rect 1490 41616 1500 41626
rect 1490 41610 1619 41616
rect 219 41576 231 41610
rect 1607 41576 1619 41610
rect 219 41570 980 41576
rect 970 41560 980 41570
rect 1490 41570 1619 41576
rect 1490 41560 1500 41570
rect 1660 41562 1706 41720
rect 342 41520 352 41530
rect 219 41514 352 41520
rect 858 41520 868 41530
rect 1660 41528 1666 41562
rect 1700 41528 1706 41562
rect 858 41514 1619 41520
rect 219 41480 231 41514
rect 1607 41480 1619 41514
rect 219 41474 352 41480
rect 132 41432 138 41466
rect 172 41432 178 41466
rect 342 41464 352 41474
rect 858 41474 1619 41480
rect 858 41464 868 41474
rect 132 41274 178 41432
rect 970 41424 980 41434
rect 219 41418 980 41424
rect 1490 41424 1500 41434
rect 1490 41418 1619 41424
rect 219 41384 231 41418
rect 1607 41384 1619 41418
rect 219 41378 980 41384
rect 970 41368 980 41378
rect 1490 41378 1619 41384
rect 1490 41368 1500 41378
rect 1660 41370 1706 41528
rect 342 41328 352 41338
rect 219 41322 352 41328
rect 858 41328 868 41338
rect 1660 41336 1666 41370
rect 1700 41336 1706 41370
rect 858 41322 1619 41328
rect 219 41288 231 41322
rect 1607 41288 1619 41322
rect 219 41282 352 41288
rect 132 41240 138 41274
rect 172 41240 178 41274
rect 342 41272 352 41282
rect 858 41282 1619 41288
rect 858 41272 868 41282
rect 132 41082 178 41240
rect 970 41232 980 41242
rect 219 41226 980 41232
rect 1490 41232 1500 41242
rect 1490 41226 1619 41232
rect 219 41192 231 41226
rect 1607 41192 1619 41226
rect 219 41186 980 41192
rect 970 41176 980 41186
rect 1490 41186 1619 41192
rect 1490 41176 1500 41186
rect 1660 41178 1706 41336
rect 342 41136 352 41146
rect 219 41130 352 41136
rect 858 41136 868 41146
rect 1660 41144 1666 41178
rect 1700 41144 1706 41178
rect 858 41130 1619 41136
rect 219 41096 231 41130
rect 1607 41096 1619 41130
rect 219 41090 352 41096
rect 132 41048 138 41082
rect 172 41048 178 41082
rect 342 41080 352 41090
rect 858 41090 1619 41096
rect 858 41080 868 41090
rect 132 40890 178 41048
rect 970 41040 980 41050
rect 219 41034 980 41040
rect 1490 41040 1500 41050
rect 1490 41034 1619 41040
rect 219 41000 231 41034
rect 1607 41000 1619 41034
rect 219 40994 980 41000
rect 970 40984 980 40994
rect 1490 40994 1619 41000
rect 1490 40984 1500 40994
rect 1660 40986 1706 41144
rect 342 40944 352 40954
rect 219 40938 352 40944
rect 858 40944 868 40954
rect 1660 40952 1666 40986
rect 1700 40952 1706 40986
rect 858 40938 1619 40944
rect 219 40904 231 40938
rect 1607 40904 1619 40938
rect 219 40898 352 40904
rect 132 40856 138 40890
rect 172 40856 178 40890
rect 342 40888 352 40898
rect 858 40898 1619 40904
rect 858 40888 868 40898
rect 132 40698 178 40856
rect 970 40848 980 40858
rect 219 40842 980 40848
rect 1490 40848 1500 40858
rect 1490 40842 1619 40848
rect 219 40808 231 40842
rect 1607 40808 1619 40842
rect 219 40802 980 40808
rect 970 40792 980 40802
rect 1490 40802 1619 40808
rect 1490 40792 1500 40802
rect 1660 40794 1706 40952
rect 342 40752 352 40762
rect 219 40746 352 40752
rect 858 40752 868 40762
rect 1660 40760 1666 40794
rect 1700 40760 1706 40794
rect 858 40746 1619 40752
rect 219 40712 231 40746
rect 1607 40712 1619 40746
rect 219 40706 352 40712
rect 132 40664 138 40698
rect 172 40664 178 40698
rect 342 40696 352 40706
rect 858 40706 1619 40712
rect 858 40696 868 40706
rect 132 40506 178 40664
rect 970 40656 980 40666
rect 219 40650 980 40656
rect 1490 40656 1500 40666
rect 1490 40650 1619 40656
rect 219 40616 231 40650
rect 1607 40616 1619 40650
rect 219 40610 980 40616
rect 970 40600 980 40610
rect 1490 40610 1619 40616
rect 1490 40600 1500 40610
rect 1660 40602 1706 40760
rect 342 40560 352 40570
rect 219 40554 352 40560
rect 858 40560 868 40570
rect 1660 40568 1666 40602
rect 1700 40568 1706 40602
rect 858 40554 1619 40560
rect 219 40520 231 40554
rect 1607 40520 1619 40554
rect 219 40514 352 40520
rect 132 40472 138 40506
rect 172 40472 178 40506
rect 342 40504 352 40514
rect 858 40514 1619 40520
rect 858 40504 868 40514
rect 132 40314 178 40472
rect 970 40464 980 40474
rect 219 40458 980 40464
rect 1490 40464 1500 40474
rect 1490 40458 1619 40464
rect 219 40424 231 40458
rect 1607 40424 1619 40458
rect 219 40418 980 40424
rect 970 40408 980 40418
rect 1490 40418 1619 40424
rect 1490 40408 1500 40418
rect 1660 40410 1706 40568
rect 342 40368 352 40378
rect 219 40362 352 40368
rect 858 40368 868 40378
rect 1660 40376 1666 40410
rect 1700 40376 1706 40410
rect 858 40362 1619 40368
rect 219 40328 231 40362
rect 1607 40328 1619 40362
rect 219 40322 352 40328
rect 132 40280 138 40314
rect 172 40280 178 40314
rect 342 40312 352 40322
rect 858 40322 1619 40328
rect 858 40312 868 40322
rect 132 40122 178 40280
rect 970 40272 980 40282
rect 219 40266 980 40272
rect 1490 40272 1500 40282
rect 1490 40266 1619 40272
rect 219 40232 231 40266
rect 1607 40232 1619 40266
rect 219 40226 980 40232
rect 970 40216 980 40226
rect 1490 40226 1619 40232
rect 1490 40216 1500 40226
rect 1660 40218 1706 40376
rect 342 40176 352 40186
rect 219 40170 352 40176
rect 858 40176 868 40186
rect 1660 40184 1666 40218
rect 1700 40184 1706 40218
rect 858 40170 1619 40176
rect 219 40136 231 40170
rect 1607 40136 1619 40170
rect 219 40130 352 40136
rect 132 40088 138 40122
rect 172 40088 178 40122
rect 342 40120 352 40130
rect 858 40130 1619 40136
rect 858 40120 868 40130
rect 132 39930 178 40088
rect 970 40080 980 40090
rect 219 40074 980 40080
rect 1490 40080 1500 40090
rect 1490 40074 1619 40080
rect 219 40040 231 40074
rect 1607 40040 1619 40074
rect 219 40034 980 40040
rect 970 40024 980 40034
rect 1490 40034 1619 40040
rect 1490 40024 1500 40034
rect 1660 40026 1706 40184
rect 342 39984 352 39994
rect 219 39978 352 39984
rect 858 39984 868 39994
rect 1660 39992 1666 40026
rect 1700 39992 1706 40026
rect 858 39978 1619 39984
rect 219 39944 231 39978
rect 1607 39944 1619 39978
rect 219 39938 352 39944
rect 132 39896 138 39930
rect 172 39896 178 39930
rect 342 39928 352 39938
rect 858 39938 1619 39944
rect 858 39928 868 39938
rect 132 39738 178 39896
rect 970 39888 980 39898
rect 219 39882 980 39888
rect 1490 39888 1500 39898
rect 1490 39882 1619 39888
rect 219 39848 231 39882
rect 1607 39848 1619 39882
rect 219 39842 980 39848
rect 970 39832 980 39842
rect 1490 39842 1619 39848
rect 1490 39832 1500 39842
rect 1660 39834 1706 39992
rect 342 39792 352 39802
rect 219 39786 352 39792
rect 858 39792 868 39802
rect 1660 39800 1666 39834
rect 1700 39800 1706 39834
rect 858 39786 1619 39792
rect 219 39752 231 39786
rect 1607 39752 1619 39786
rect 219 39746 352 39752
rect 132 39704 138 39738
rect 172 39704 178 39738
rect 342 39736 352 39746
rect 858 39746 1619 39752
rect 858 39736 868 39746
rect 132 39546 178 39704
rect 970 39696 980 39706
rect 219 39690 980 39696
rect 1490 39696 1500 39706
rect 1490 39690 1619 39696
rect 219 39656 231 39690
rect 1607 39656 1619 39690
rect 219 39650 980 39656
rect 970 39640 980 39650
rect 1490 39650 1619 39656
rect 1490 39640 1500 39650
rect 1660 39642 1706 39800
rect 342 39600 352 39610
rect 219 39594 352 39600
rect 858 39600 868 39610
rect 1660 39608 1666 39642
rect 1700 39608 1706 39642
rect 858 39594 1619 39600
rect 219 39560 231 39594
rect 1607 39560 1619 39594
rect 219 39554 352 39560
rect 132 39512 138 39546
rect 172 39512 178 39546
rect 342 39544 352 39554
rect 858 39554 1619 39560
rect 858 39544 868 39554
rect 132 39354 178 39512
rect 970 39504 980 39514
rect 219 39498 980 39504
rect 1490 39504 1500 39514
rect 1490 39498 1619 39504
rect 219 39464 231 39498
rect 1607 39464 1619 39498
rect 219 39458 980 39464
rect 970 39448 980 39458
rect 1490 39458 1619 39464
rect 1490 39448 1500 39458
rect 1660 39450 1706 39608
rect 342 39408 352 39418
rect 219 39402 352 39408
rect 858 39408 868 39418
rect 1660 39416 1666 39450
rect 1700 39416 1706 39450
rect 858 39402 1619 39408
rect 219 39368 231 39402
rect 1607 39368 1619 39402
rect 219 39362 352 39368
rect 132 39320 138 39354
rect 172 39320 178 39354
rect 342 39352 352 39362
rect 858 39362 1619 39368
rect 858 39352 868 39362
rect 132 39162 178 39320
rect 970 39312 980 39322
rect 219 39306 980 39312
rect 1490 39312 1500 39322
rect 1490 39306 1619 39312
rect 219 39272 231 39306
rect 1607 39272 1619 39306
rect 219 39266 980 39272
rect 970 39256 980 39266
rect 1490 39266 1619 39272
rect 1490 39256 1500 39266
rect 1660 39258 1706 39416
rect 342 39216 352 39226
rect 219 39210 352 39216
rect 858 39216 868 39226
rect 1660 39224 1666 39258
rect 1700 39224 1706 39258
rect 858 39210 1619 39216
rect 219 39176 231 39210
rect 1607 39176 1619 39210
rect 219 39170 352 39176
rect 132 39128 138 39162
rect 172 39128 178 39162
rect 342 39160 352 39170
rect 858 39170 1619 39176
rect 858 39160 868 39170
rect 132 38970 178 39128
rect 970 39120 980 39130
rect 219 39114 980 39120
rect 1490 39120 1500 39130
rect 1490 39114 1619 39120
rect 219 39080 231 39114
rect 1607 39080 1619 39114
rect 219 39074 980 39080
rect 970 39064 980 39074
rect 1490 39074 1619 39080
rect 1490 39064 1500 39074
rect 1660 39066 1706 39224
rect 342 39024 352 39034
rect 219 39018 352 39024
rect 858 39024 868 39034
rect 1660 39032 1666 39066
rect 1700 39032 1706 39066
rect 858 39018 1619 39024
rect 219 38984 231 39018
rect 1607 38984 1619 39018
rect 219 38978 352 38984
rect 132 38936 138 38970
rect 172 38936 178 38970
rect 342 38968 352 38978
rect 858 38978 1619 38984
rect 858 38968 868 38978
rect 132 38778 178 38936
rect 970 38928 980 38938
rect 219 38922 980 38928
rect 1490 38928 1500 38938
rect 1490 38922 1619 38928
rect 219 38888 231 38922
rect 1607 38888 1619 38922
rect 219 38882 980 38888
rect 970 38872 980 38882
rect 1490 38882 1619 38888
rect 1490 38872 1500 38882
rect 1660 38874 1706 39032
rect 342 38832 352 38842
rect 219 38826 352 38832
rect 858 38832 868 38842
rect 1660 38840 1666 38874
rect 1700 38840 1706 38874
rect 858 38826 1619 38832
rect 219 38792 231 38826
rect 1607 38792 1619 38826
rect 219 38786 352 38792
rect 132 38744 138 38778
rect 172 38744 178 38778
rect 342 38776 352 38786
rect 858 38786 1619 38792
rect 858 38776 868 38786
rect 132 38586 178 38744
rect 970 38736 980 38746
rect 219 38730 980 38736
rect 1490 38736 1500 38746
rect 1490 38730 1619 38736
rect 219 38696 231 38730
rect 1607 38696 1619 38730
rect 219 38690 980 38696
rect 970 38680 980 38690
rect 1490 38690 1619 38696
rect 1490 38680 1500 38690
rect 1660 38682 1706 38840
rect 342 38640 352 38650
rect 219 38634 352 38640
rect 858 38640 868 38650
rect 1660 38648 1666 38682
rect 1700 38648 1706 38682
rect 858 38634 1619 38640
rect 219 38600 231 38634
rect 1607 38600 1619 38634
rect 219 38594 352 38600
rect 132 38552 138 38586
rect 172 38552 178 38586
rect 342 38584 352 38594
rect 858 38594 1619 38600
rect 858 38584 868 38594
rect 132 38394 178 38552
rect 970 38544 980 38554
rect 219 38538 980 38544
rect 1490 38544 1500 38554
rect 1490 38538 1619 38544
rect 219 38504 231 38538
rect 1607 38504 1619 38538
rect 219 38498 980 38504
rect 970 38488 980 38498
rect 1490 38498 1619 38504
rect 1490 38488 1500 38498
rect 1660 38490 1706 38648
rect 342 38448 352 38458
rect 219 38442 352 38448
rect 858 38448 868 38458
rect 1660 38456 1666 38490
rect 1700 38456 1706 38490
rect 858 38442 1619 38448
rect 219 38408 231 38442
rect 1607 38408 1619 38442
rect 219 38402 352 38408
rect 132 38360 138 38394
rect 172 38360 178 38394
rect 342 38392 352 38402
rect 858 38402 1619 38408
rect 858 38392 868 38402
rect 132 38202 178 38360
rect 970 38352 980 38362
rect 219 38346 980 38352
rect 1490 38352 1500 38362
rect 1490 38346 1619 38352
rect 219 38312 231 38346
rect 1607 38312 1619 38346
rect 219 38306 980 38312
rect 970 38296 980 38306
rect 1490 38306 1619 38312
rect 1490 38296 1500 38306
rect 1660 38298 1706 38456
rect 342 38256 352 38266
rect 219 38250 352 38256
rect 858 38256 868 38266
rect 1660 38264 1666 38298
rect 1700 38264 1706 38298
rect 858 38250 1619 38256
rect 219 38216 231 38250
rect 1607 38216 1619 38250
rect 219 38210 352 38216
rect 132 38168 138 38202
rect 172 38168 178 38202
rect 342 38200 352 38210
rect 858 38210 1619 38216
rect 858 38200 868 38210
rect 132 38010 178 38168
rect 970 38160 980 38170
rect 219 38154 980 38160
rect 1490 38160 1500 38170
rect 1490 38154 1619 38160
rect 219 38120 231 38154
rect 1607 38120 1619 38154
rect 219 38114 980 38120
rect 970 38104 980 38114
rect 1490 38114 1619 38120
rect 1490 38104 1500 38114
rect 1660 38106 1706 38264
rect 342 38064 352 38074
rect 219 38058 352 38064
rect 858 38064 868 38074
rect 1660 38072 1666 38106
rect 1700 38072 1706 38106
rect 858 38058 1619 38064
rect 219 38024 231 38058
rect 1607 38024 1619 38058
rect 219 38018 352 38024
rect 132 37976 138 38010
rect 172 37976 178 38010
rect 342 38008 352 38018
rect 858 38018 1619 38024
rect 858 38008 868 38018
rect 132 37818 178 37976
rect 970 37968 980 37978
rect 219 37962 980 37968
rect 1490 37968 1500 37978
rect 1490 37962 1619 37968
rect 219 37928 231 37962
rect 1607 37928 1619 37962
rect 219 37922 980 37928
rect 970 37912 980 37922
rect 1490 37922 1619 37928
rect 1490 37912 1500 37922
rect 1660 37914 1706 38072
rect 342 37872 352 37882
rect 219 37866 352 37872
rect 858 37872 868 37882
rect 1660 37880 1666 37914
rect 1700 37880 1706 37914
rect 858 37866 1619 37872
rect 219 37832 231 37866
rect 1607 37832 1619 37866
rect 219 37826 352 37832
rect 132 37784 138 37818
rect 172 37784 178 37818
rect 342 37816 352 37826
rect 858 37826 1619 37832
rect 858 37816 868 37826
rect 132 37626 178 37784
rect 970 37776 980 37786
rect 219 37770 980 37776
rect 1490 37776 1500 37786
rect 1490 37770 1619 37776
rect 219 37736 231 37770
rect 1607 37736 1619 37770
rect 219 37730 980 37736
rect 970 37720 980 37730
rect 1490 37730 1619 37736
rect 1490 37720 1500 37730
rect 1660 37722 1706 37880
rect 342 37680 352 37690
rect 219 37674 352 37680
rect 858 37680 868 37690
rect 1660 37688 1666 37722
rect 1700 37688 1706 37722
rect 858 37674 1619 37680
rect 219 37640 231 37674
rect 1607 37640 1619 37674
rect 219 37634 352 37640
rect 132 37592 138 37626
rect 172 37592 178 37626
rect 342 37624 352 37634
rect 858 37634 1619 37640
rect 858 37624 868 37634
rect 132 37434 178 37592
rect 970 37584 980 37594
rect 219 37578 980 37584
rect 1490 37584 1500 37594
rect 1490 37578 1619 37584
rect 219 37544 231 37578
rect 1607 37544 1619 37578
rect 219 37538 980 37544
rect 970 37528 980 37538
rect 1490 37538 1619 37544
rect 1490 37528 1500 37538
rect 1660 37530 1706 37688
rect 342 37488 352 37498
rect 219 37482 352 37488
rect 858 37488 868 37498
rect 1660 37496 1666 37530
rect 1700 37496 1706 37530
rect 858 37482 1619 37488
rect 219 37448 231 37482
rect 1607 37448 1619 37482
rect 219 37442 352 37448
rect 132 37400 138 37434
rect 172 37400 178 37434
rect 342 37432 352 37442
rect 858 37442 1619 37448
rect 858 37432 868 37442
rect 132 37242 178 37400
rect 970 37392 980 37402
rect 219 37386 980 37392
rect 1490 37392 1500 37402
rect 1490 37386 1619 37392
rect 219 37352 231 37386
rect 1607 37352 1619 37386
rect 219 37346 980 37352
rect 970 37336 980 37346
rect 1490 37346 1619 37352
rect 1490 37336 1500 37346
rect 1660 37338 1706 37496
rect 342 37296 352 37306
rect 219 37290 352 37296
rect 858 37296 868 37306
rect 1660 37304 1666 37338
rect 1700 37304 1706 37338
rect 858 37290 1619 37296
rect 219 37256 231 37290
rect 1607 37256 1619 37290
rect 219 37250 352 37256
rect 132 37208 138 37242
rect 172 37208 178 37242
rect 342 37240 352 37250
rect 858 37250 1619 37256
rect 858 37240 868 37250
rect 132 37050 178 37208
rect 970 37200 980 37210
rect 219 37194 980 37200
rect 1490 37200 1500 37210
rect 1490 37194 1619 37200
rect 219 37160 231 37194
rect 1607 37160 1619 37194
rect 219 37154 980 37160
rect 970 37144 980 37154
rect 1490 37154 1619 37160
rect 1490 37144 1500 37154
rect 1660 37146 1706 37304
rect 342 37104 352 37114
rect 219 37098 352 37104
rect 858 37104 868 37114
rect 1660 37112 1666 37146
rect 1700 37112 1706 37146
rect 858 37098 1619 37104
rect 219 37064 231 37098
rect 1607 37064 1619 37098
rect 219 37058 352 37064
rect 132 37016 138 37050
rect 172 37016 178 37050
rect 342 37048 352 37058
rect 858 37058 1619 37064
rect 858 37048 868 37058
rect 132 36858 178 37016
rect 970 37008 980 37018
rect 219 37002 980 37008
rect 1490 37008 1500 37018
rect 1490 37002 1619 37008
rect 219 36968 231 37002
rect 1607 36968 1619 37002
rect 219 36962 980 36968
rect 970 36952 980 36962
rect 1490 36962 1619 36968
rect 1490 36952 1500 36962
rect 1660 36954 1706 37112
rect 342 36912 352 36922
rect 219 36906 352 36912
rect 858 36912 868 36922
rect 1660 36920 1666 36954
rect 1700 36920 1706 36954
rect 858 36906 1619 36912
rect 219 36872 231 36906
rect 1607 36872 1619 36906
rect 219 36866 352 36872
rect 132 36824 138 36858
rect 172 36824 178 36858
rect 342 36856 352 36866
rect 858 36866 1619 36872
rect 858 36856 868 36866
rect 132 36666 178 36824
rect 970 36816 980 36826
rect 219 36810 980 36816
rect 1490 36816 1500 36826
rect 1490 36810 1619 36816
rect 219 36776 231 36810
rect 1607 36776 1619 36810
rect 219 36770 980 36776
rect 970 36760 980 36770
rect 1490 36770 1619 36776
rect 1490 36760 1500 36770
rect 1660 36762 1706 36920
rect 342 36720 352 36730
rect 219 36714 352 36720
rect 858 36720 868 36730
rect 1660 36728 1666 36762
rect 1700 36728 1706 36762
rect 858 36714 1619 36720
rect 219 36680 231 36714
rect 1607 36680 1619 36714
rect 219 36674 352 36680
rect 132 36632 138 36666
rect 172 36632 178 36666
rect 342 36664 352 36674
rect 858 36674 1619 36680
rect 858 36664 868 36674
rect 132 36474 178 36632
rect 970 36624 980 36634
rect 219 36618 980 36624
rect 1490 36624 1500 36634
rect 1490 36618 1619 36624
rect 219 36584 231 36618
rect 1607 36584 1619 36618
rect 219 36578 980 36584
rect 970 36568 980 36578
rect 1490 36578 1619 36584
rect 1490 36568 1500 36578
rect 1660 36570 1706 36728
rect 342 36528 352 36538
rect 219 36522 352 36528
rect 858 36528 868 36538
rect 1660 36536 1666 36570
rect 1700 36536 1706 36570
rect 858 36522 1619 36528
rect 219 36488 231 36522
rect 1607 36488 1619 36522
rect 219 36482 352 36488
rect 132 36440 138 36474
rect 172 36440 178 36474
rect 342 36472 352 36482
rect 858 36482 1619 36488
rect 858 36472 868 36482
rect 132 36282 178 36440
rect 970 36432 980 36442
rect 219 36426 980 36432
rect 1490 36432 1500 36442
rect 1490 36426 1619 36432
rect 219 36392 231 36426
rect 1607 36392 1619 36426
rect 219 36386 980 36392
rect 970 36376 980 36386
rect 1490 36386 1619 36392
rect 1490 36376 1500 36386
rect 1660 36378 1706 36536
rect 342 36336 352 36346
rect 219 36330 352 36336
rect 858 36336 868 36346
rect 1660 36344 1666 36378
rect 1700 36344 1706 36378
rect 858 36330 1619 36336
rect 219 36296 231 36330
rect 1607 36296 1619 36330
rect 219 36290 352 36296
rect 132 36248 138 36282
rect 172 36248 178 36282
rect 342 36280 352 36290
rect 858 36290 1619 36296
rect 858 36280 868 36290
rect 132 36090 178 36248
rect 970 36240 980 36250
rect 219 36234 980 36240
rect 1490 36240 1500 36250
rect 1490 36234 1619 36240
rect 219 36200 231 36234
rect 1607 36200 1619 36234
rect 219 36194 980 36200
rect 970 36184 980 36194
rect 1490 36194 1619 36200
rect 1490 36184 1500 36194
rect 1660 36186 1706 36344
rect 342 36144 352 36154
rect 219 36138 352 36144
rect 858 36144 868 36154
rect 1660 36152 1666 36186
rect 1700 36152 1706 36186
rect 858 36138 1619 36144
rect 219 36104 231 36138
rect 1607 36104 1619 36138
rect 219 36098 352 36104
rect 132 36056 138 36090
rect 172 36056 178 36090
rect 342 36088 352 36098
rect 858 36098 1619 36104
rect 858 36088 868 36098
rect 132 35898 178 36056
rect 970 36048 980 36058
rect 219 36042 980 36048
rect 1490 36048 1500 36058
rect 1490 36042 1619 36048
rect 219 36008 231 36042
rect 1607 36008 1619 36042
rect 219 36002 980 36008
rect 970 35992 980 36002
rect 1490 36002 1619 36008
rect 1490 35992 1500 36002
rect 1660 35994 1706 36152
rect 342 35952 352 35962
rect 219 35946 352 35952
rect 858 35952 868 35962
rect 1660 35960 1666 35994
rect 1700 35960 1706 35994
rect 858 35946 1619 35952
rect 219 35912 231 35946
rect 1607 35912 1619 35946
rect 219 35906 352 35912
rect 132 35864 138 35898
rect 172 35864 178 35898
rect 342 35896 352 35906
rect 858 35906 1619 35912
rect 858 35896 868 35906
rect 132 35706 178 35864
rect 970 35856 980 35866
rect 219 35850 980 35856
rect 1490 35856 1500 35866
rect 1490 35850 1619 35856
rect 219 35816 231 35850
rect 1607 35816 1619 35850
rect 219 35810 980 35816
rect 970 35800 980 35810
rect 1490 35810 1619 35816
rect 1490 35800 1500 35810
rect 1660 35802 1706 35960
rect 342 35760 352 35770
rect 219 35754 352 35760
rect 858 35760 868 35770
rect 1660 35768 1666 35802
rect 1700 35768 1706 35802
rect 858 35754 1619 35760
rect 219 35720 231 35754
rect 1607 35720 1619 35754
rect 219 35714 352 35720
rect 132 35672 138 35706
rect 172 35672 178 35706
rect 342 35704 352 35714
rect 858 35714 1619 35720
rect 858 35704 868 35714
rect 132 35514 178 35672
rect 970 35664 980 35674
rect 219 35658 980 35664
rect 1490 35664 1500 35674
rect 1490 35658 1619 35664
rect 219 35624 231 35658
rect 1607 35624 1619 35658
rect 219 35618 980 35624
rect 970 35608 980 35618
rect 1490 35618 1619 35624
rect 1490 35608 1500 35618
rect 1660 35610 1706 35768
rect 342 35568 352 35578
rect 219 35562 352 35568
rect 858 35568 868 35578
rect 1660 35576 1666 35610
rect 1700 35576 1706 35610
rect 858 35562 1619 35568
rect 219 35528 231 35562
rect 1607 35528 1619 35562
rect 219 35522 352 35528
rect 132 35480 138 35514
rect 172 35480 178 35514
rect 342 35512 352 35522
rect 858 35522 1619 35528
rect 858 35512 868 35522
rect 132 35322 178 35480
rect 970 35472 980 35482
rect 219 35466 980 35472
rect 1490 35472 1500 35482
rect 1490 35466 1619 35472
rect 219 35432 231 35466
rect 1607 35432 1619 35466
rect 219 35426 980 35432
rect 970 35416 980 35426
rect 1490 35426 1619 35432
rect 1490 35416 1500 35426
rect 1660 35418 1706 35576
rect 342 35376 352 35386
rect 219 35370 352 35376
rect 858 35376 868 35386
rect 1660 35384 1666 35418
rect 1700 35384 1706 35418
rect 858 35370 1619 35376
rect 219 35336 231 35370
rect 1607 35336 1619 35370
rect 219 35330 352 35336
rect 132 35288 138 35322
rect 172 35288 178 35322
rect 342 35320 352 35330
rect 858 35330 1619 35336
rect 858 35320 868 35330
rect 132 35130 178 35288
rect 970 35280 980 35290
rect 219 35274 980 35280
rect 1490 35280 1500 35290
rect 1490 35274 1619 35280
rect 219 35240 231 35274
rect 1607 35240 1619 35274
rect 219 35234 980 35240
rect 970 35224 980 35234
rect 1490 35234 1619 35240
rect 1490 35224 1500 35234
rect 1660 35226 1706 35384
rect 342 35184 352 35194
rect 219 35178 352 35184
rect 858 35184 868 35194
rect 1660 35192 1666 35226
rect 1700 35192 1706 35226
rect 858 35178 1619 35184
rect 219 35144 231 35178
rect 1607 35144 1619 35178
rect 219 35138 352 35144
rect 132 35096 138 35130
rect 172 35096 178 35130
rect 342 35128 352 35138
rect 858 35138 1619 35144
rect 858 35128 868 35138
rect 132 34938 178 35096
rect 970 35088 980 35098
rect 219 35082 980 35088
rect 1490 35088 1500 35098
rect 1490 35082 1619 35088
rect 219 35048 231 35082
rect 1607 35048 1619 35082
rect 219 35042 980 35048
rect 970 35032 980 35042
rect 1490 35042 1619 35048
rect 1490 35032 1500 35042
rect 1660 35034 1706 35192
rect 342 34992 352 35002
rect 219 34986 352 34992
rect 858 34992 868 35002
rect 1660 35000 1666 35034
rect 1700 35000 1706 35034
rect 858 34986 1619 34992
rect 219 34952 231 34986
rect 1607 34952 1619 34986
rect 219 34946 352 34952
rect 132 34904 138 34938
rect 172 34904 178 34938
rect 342 34936 352 34946
rect 858 34946 1619 34952
rect 858 34936 868 34946
rect 132 34746 178 34904
rect 970 34896 980 34906
rect 219 34890 980 34896
rect 1490 34896 1500 34906
rect 1490 34890 1619 34896
rect 219 34856 231 34890
rect 1607 34856 1619 34890
rect 219 34850 980 34856
rect 970 34840 980 34850
rect 1490 34850 1619 34856
rect 1490 34840 1500 34850
rect 1660 34842 1706 35000
rect 342 34800 352 34810
rect 219 34794 352 34800
rect 858 34800 868 34810
rect 1660 34808 1666 34842
rect 1700 34808 1706 34842
rect 858 34794 1619 34800
rect 219 34760 231 34794
rect 1607 34760 1619 34794
rect 219 34754 352 34760
rect 132 34712 138 34746
rect 172 34712 178 34746
rect 342 34744 352 34754
rect 858 34754 1619 34760
rect 858 34744 868 34754
rect 132 34554 178 34712
rect 970 34704 980 34714
rect 219 34698 980 34704
rect 1490 34704 1500 34714
rect 1490 34698 1619 34704
rect 219 34664 231 34698
rect 1607 34664 1619 34698
rect 219 34658 980 34664
rect 970 34648 980 34658
rect 1490 34658 1619 34664
rect 1490 34648 1500 34658
rect 1660 34650 1706 34808
rect 342 34608 352 34618
rect 219 34602 352 34608
rect 858 34608 868 34618
rect 1660 34616 1666 34650
rect 1700 34616 1706 34650
rect 858 34602 1619 34608
rect 219 34568 231 34602
rect 1607 34568 1619 34602
rect 219 34562 352 34568
rect 132 34520 138 34554
rect 172 34520 178 34554
rect 342 34552 352 34562
rect 858 34562 1619 34568
rect 858 34552 868 34562
rect 132 34362 178 34520
rect 970 34512 980 34522
rect 219 34506 980 34512
rect 1490 34512 1500 34522
rect 1490 34506 1619 34512
rect 219 34472 231 34506
rect 1607 34472 1619 34506
rect 219 34466 980 34472
rect 970 34456 980 34466
rect 1490 34466 1619 34472
rect 1490 34456 1500 34466
rect 1660 34458 1706 34616
rect 342 34416 352 34426
rect 219 34410 352 34416
rect 858 34416 868 34426
rect 1660 34424 1666 34458
rect 1700 34424 1706 34458
rect 858 34410 1619 34416
rect 219 34376 231 34410
rect 1607 34376 1619 34410
rect 219 34370 352 34376
rect 132 34328 138 34362
rect 172 34328 178 34362
rect 342 34360 352 34370
rect 858 34370 1619 34376
rect 858 34360 868 34370
rect 132 34170 178 34328
rect 970 34320 980 34330
rect 219 34314 980 34320
rect 1490 34320 1500 34330
rect 1490 34314 1619 34320
rect 219 34280 231 34314
rect 1607 34280 1619 34314
rect 219 34274 980 34280
rect 970 34264 980 34274
rect 1490 34274 1619 34280
rect 1490 34264 1500 34274
rect 1660 34266 1706 34424
rect 342 34224 352 34234
rect 219 34218 352 34224
rect 858 34224 868 34234
rect 1660 34232 1666 34266
rect 1700 34232 1706 34266
rect 858 34218 1619 34224
rect 219 34184 231 34218
rect 1607 34184 1619 34218
rect 219 34178 352 34184
rect 132 34136 138 34170
rect 172 34136 178 34170
rect 342 34168 352 34178
rect 858 34178 1619 34184
rect 858 34168 868 34178
rect 132 33978 178 34136
rect 970 34128 980 34138
rect 219 34122 980 34128
rect 1490 34128 1500 34138
rect 1490 34122 1619 34128
rect 219 34088 231 34122
rect 1607 34088 1619 34122
rect 219 34082 980 34088
rect 970 34072 980 34082
rect 1490 34082 1619 34088
rect 1490 34072 1500 34082
rect 1660 34074 1706 34232
rect 342 34032 352 34042
rect 219 34026 352 34032
rect 858 34032 868 34042
rect 1660 34040 1666 34074
rect 1700 34040 1706 34074
rect 858 34026 1619 34032
rect 219 33992 231 34026
rect 1607 33992 1619 34026
rect 219 33986 352 33992
rect 132 33944 138 33978
rect 172 33944 178 33978
rect 342 33976 352 33986
rect 858 33986 1619 33992
rect 858 33976 868 33986
rect 132 33786 178 33944
rect 970 33936 980 33946
rect 219 33930 980 33936
rect 1490 33936 1500 33946
rect 1490 33930 1619 33936
rect 219 33896 231 33930
rect 1607 33896 1619 33930
rect 219 33890 980 33896
rect 970 33880 980 33890
rect 1490 33890 1619 33896
rect 1490 33880 1500 33890
rect 1660 33882 1706 34040
rect 342 33840 352 33850
rect 219 33834 352 33840
rect 858 33840 868 33850
rect 1660 33848 1666 33882
rect 1700 33848 1706 33882
rect 858 33834 1619 33840
rect 219 33800 231 33834
rect 1607 33800 1619 33834
rect 219 33794 352 33800
rect 132 33752 138 33786
rect 172 33752 178 33786
rect 342 33784 352 33794
rect 858 33794 1619 33800
rect 858 33784 868 33794
rect 132 33594 178 33752
rect 970 33744 980 33754
rect 219 33738 980 33744
rect 1490 33744 1500 33754
rect 1490 33738 1619 33744
rect 219 33704 231 33738
rect 1607 33704 1619 33738
rect 219 33698 980 33704
rect 970 33688 980 33698
rect 1490 33698 1619 33704
rect 1490 33688 1500 33698
rect 1660 33690 1706 33848
rect 342 33648 352 33658
rect 219 33642 352 33648
rect 858 33648 868 33658
rect 1660 33656 1666 33690
rect 1700 33656 1706 33690
rect 858 33642 1619 33648
rect 219 33608 231 33642
rect 1607 33608 1619 33642
rect 219 33602 352 33608
rect 132 33560 138 33594
rect 172 33560 178 33594
rect 342 33592 352 33602
rect 858 33602 1619 33608
rect 858 33592 868 33602
rect 132 33402 178 33560
rect 970 33552 980 33562
rect 219 33546 980 33552
rect 1490 33552 1500 33562
rect 1490 33546 1619 33552
rect 219 33512 231 33546
rect 1607 33512 1619 33546
rect 219 33506 980 33512
rect 970 33496 980 33506
rect 1490 33506 1619 33512
rect 1490 33496 1500 33506
rect 1660 33498 1706 33656
rect 342 33456 352 33466
rect 219 33450 352 33456
rect 858 33456 868 33466
rect 1660 33464 1666 33498
rect 1700 33464 1706 33498
rect 858 33450 1619 33456
rect 219 33416 231 33450
rect 1607 33416 1619 33450
rect 219 33410 352 33416
rect 132 33368 138 33402
rect 172 33368 178 33402
rect 342 33400 352 33410
rect 858 33410 1619 33416
rect 858 33400 868 33410
rect 132 33210 178 33368
rect 970 33360 980 33370
rect 219 33354 980 33360
rect 1490 33360 1500 33370
rect 1490 33354 1619 33360
rect 219 33320 231 33354
rect 1607 33320 1619 33354
rect 219 33314 980 33320
rect 970 33304 980 33314
rect 1490 33314 1619 33320
rect 1490 33304 1500 33314
rect 1660 33306 1706 33464
rect 342 33264 352 33274
rect 219 33258 352 33264
rect 858 33264 868 33274
rect 1660 33272 1666 33306
rect 1700 33272 1706 33306
rect 858 33258 1619 33264
rect 219 33224 231 33258
rect 1607 33224 1619 33258
rect 219 33218 352 33224
rect 132 33176 138 33210
rect 172 33176 178 33210
rect 342 33208 352 33218
rect 858 33218 1619 33224
rect 858 33208 868 33218
rect 132 33018 178 33176
rect 970 33168 980 33178
rect 219 33162 980 33168
rect 1490 33168 1500 33178
rect 1490 33162 1619 33168
rect 219 33128 231 33162
rect 1607 33128 1619 33162
rect 219 33122 980 33128
rect 970 33112 980 33122
rect 1490 33122 1619 33128
rect 1490 33112 1500 33122
rect 1660 33114 1706 33272
rect 342 33072 352 33082
rect 219 33066 352 33072
rect 858 33072 868 33082
rect 1660 33080 1666 33114
rect 1700 33080 1706 33114
rect 858 33066 1619 33072
rect 219 33032 231 33066
rect 1607 33032 1619 33066
rect 219 33026 352 33032
rect 132 32984 138 33018
rect 172 32984 178 33018
rect 342 33016 352 33026
rect 858 33026 1619 33032
rect 858 33016 868 33026
rect 132 32826 178 32984
rect 970 32976 980 32986
rect 219 32970 980 32976
rect 1490 32976 1500 32986
rect 1490 32970 1619 32976
rect 219 32936 231 32970
rect 1607 32936 1619 32970
rect 219 32930 980 32936
rect 970 32920 980 32930
rect 1490 32930 1619 32936
rect 1490 32920 1500 32930
rect 1660 32922 1706 33080
rect 342 32880 352 32890
rect 219 32874 352 32880
rect 858 32880 868 32890
rect 1660 32888 1666 32922
rect 1700 32888 1706 32922
rect 858 32874 1619 32880
rect 219 32840 231 32874
rect 1607 32840 1619 32874
rect 219 32834 352 32840
rect 132 32792 138 32826
rect 172 32792 178 32826
rect 342 32824 352 32834
rect 858 32834 1619 32840
rect 858 32824 868 32834
rect 132 32634 178 32792
rect 970 32784 980 32794
rect 219 32778 980 32784
rect 1490 32784 1500 32794
rect 1490 32778 1619 32784
rect 219 32744 231 32778
rect 1607 32744 1619 32778
rect 219 32738 980 32744
rect 970 32728 980 32738
rect 1490 32738 1619 32744
rect 1490 32728 1500 32738
rect 1660 32730 1706 32888
rect 342 32688 352 32698
rect 219 32682 352 32688
rect 858 32688 868 32698
rect 1660 32696 1666 32730
rect 1700 32696 1706 32730
rect 858 32682 1619 32688
rect 219 32648 231 32682
rect 1607 32648 1619 32682
rect 219 32642 352 32648
rect 132 32600 138 32634
rect 172 32600 178 32634
rect 342 32632 352 32642
rect 858 32642 1619 32648
rect 858 32632 868 32642
rect 132 32442 178 32600
rect 970 32592 980 32602
rect 219 32586 980 32592
rect 1490 32592 1500 32602
rect 1490 32586 1619 32592
rect 219 32552 231 32586
rect 1607 32552 1619 32586
rect 219 32546 980 32552
rect 970 32536 980 32546
rect 1490 32546 1619 32552
rect 1490 32536 1500 32546
rect 1660 32538 1706 32696
rect 342 32496 352 32506
rect 219 32490 352 32496
rect 858 32496 868 32506
rect 1660 32504 1666 32538
rect 1700 32504 1706 32538
rect 858 32490 1619 32496
rect 219 32456 231 32490
rect 1607 32456 1619 32490
rect 219 32450 352 32456
rect 132 32408 138 32442
rect 172 32408 178 32442
rect 342 32440 352 32450
rect 858 32450 1619 32456
rect 858 32440 868 32450
rect 132 32250 178 32408
rect 970 32400 980 32410
rect 219 32394 980 32400
rect 1490 32400 1500 32410
rect 1490 32394 1619 32400
rect 219 32360 231 32394
rect 1607 32360 1619 32394
rect 219 32354 980 32360
rect 970 32344 980 32354
rect 1490 32354 1619 32360
rect 1490 32344 1500 32354
rect 1660 32346 1706 32504
rect 342 32304 352 32314
rect 219 32298 352 32304
rect 858 32304 868 32314
rect 1660 32312 1666 32346
rect 1700 32312 1706 32346
rect 858 32298 1619 32304
rect 219 32264 231 32298
rect 1607 32264 1619 32298
rect 219 32258 352 32264
rect 132 32216 138 32250
rect 172 32216 178 32250
rect 342 32248 352 32258
rect 858 32258 1619 32264
rect 858 32248 868 32258
rect 132 32058 178 32216
rect 970 32208 980 32218
rect 219 32202 980 32208
rect 1490 32208 1500 32218
rect 1490 32202 1619 32208
rect 219 32168 231 32202
rect 1607 32168 1619 32202
rect 219 32162 980 32168
rect 970 32152 980 32162
rect 1490 32162 1619 32168
rect 1490 32152 1500 32162
rect 1660 32154 1706 32312
rect 342 32112 352 32122
rect 219 32106 352 32112
rect 858 32112 868 32122
rect 1660 32120 1666 32154
rect 1700 32120 1706 32154
rect 858 32106 1619 32112
rect 219 32072 231 32106
rect 1607 32072 1619 32106
rect 219 32066 352 32072
rect 132 32024 138 32058
rect 172 32024 178 32058
rect 342 32056 352 32066
rect 858 32066 1619 32072
rect 858 32056 868 32066
rect 132 31866 178 32024
rect 970 32016 980 32026
rect 219 32010 980 32016
rect 1490 32016 1500 32026
rect 1490 32010 1619 32016
rect 219 31976 231 32010
rect 1607 31976 1619 32010
rect 219 31970 980 31976
rect 970 31960 980 31970
rect 1490 31970 1619 31976
rect 1490 31960 1500 31970
rect 1660 31962 1706 32120
rect 342 31920 352 31930
rect 219 31914 352 31920
rect 858 31920 868 31930
rect 1660 31928 1666 31962
rect 1700 31928 1706 31962
rect 858 31914 1619 31920
rect 219 31880 231 31914
rect 1607 31880 1619 31914
rect 219 31874 352 31880
rect 132 31832 138 31866
rect 172 31832 178 31866
rect 342 31864 352 31874
rect 858 31874 1619 31880
rect 858 31864 868 31874
rect 132 31674 178 31832
rect 970 31824 980 31834
rect 219 31818 980 31824
rect 1490 31824 1500 31834
rect 1490 31818 1619 31824
rect 219 31784 231 31818
rect 1607 31784 1619 31818
rect 219 31778 980 31784
rect 970 31768 980 31778
rect 1490 31778 1619 31784
rect 1490 31768 1500 31778
rect 1660 31770 1706 31928
rect 342 31728 352 31738
rect 219 31722 352 31728
rect 858 31728 868 31738
rect 1660 31736 1666 31770
rect 1700 31736 1706 31770
rect 858 31722 1619 31728
rect 219 31688 231 31722
rect 1607 31688 1619 31722
rect 219 31682 352 31688
rect 132 31640 138 31674
rect 172 31640 178 31674
rect 342 31672 352 31682
rect 858 31682 1619 31688
rect 858 31672 868 31682
rect 132 31482 178 31640
rect 970 31632 980 31642
rect 219 31626 980 31632
rect 1490 31632 1500 31642
rect 1490 31626 1619 31632
rect 219 31592 231 31626
rect 1607 31592 1619 31626
rect 219 31586 980 31592
rect 970 31576 980 31586
rect 1490 31586 1619 31592
rect 1490 31576 1500 31586
rect 1660 31578 1706 31736
rect 342 31536 352 31546
rect 219 31530 352 31536
rect 858 31536 868 31546
rect 1660 31544 1666 31578
rect 1700 31544 1706 31578
rect 858 31530 1619 31536
rect 219 31496 231 31530
rect 1607 31496 1619 31530
rect 219 31490 352 31496
rect 132 31448 138 31482
rect 172 31448 178 31482
rect 342 31480 352 31490
rect 858 31490 1619 31496
rect 858 31480 868 31490
rect 132 31290 178 31448
rect 970 31440 980 31450
rect 219 31434 980 31440
rect 1490 31440 1500 31450
rect 1490 31434 1619 31440
rect 219 31400 231 31434
rect 1607 31400 1619 31434
rect 219 31394 980 31400
rect 970 31384 980 31394
rect 1490 31394 1619 31400
rect 1490 31384 1500 31394
rect 1660 31386 1706 31544
rect 342 31344 352 31354
rect 219 31338 352 31344
rect 858 31344 868 31354
rect 1660 31352 1666 31386
rect 1700 31352 1706 31386
rect 858 31338 1619 31344
rect 219 31304 231 31338
rect 1607 31304 1619 31338
rect 219 31298 352 31304
rect 132 31256 138 31290
rect 172 31256 178 31290
rect 342 31288 352 31298
rect 858 31298 1619 31304
rect 858 31288 868 31298
rect 132 31098 178 31256
rect 970 31248 980 31258
rect 219 31242 980 31248
rect 1490 31248 1500 31258
rect 1490 31242 1619 31248
rect 219 31208 231 31242
rect 1607 31208 1619 31242
rect 219 31202 980 31208
rect 970 31192 980 31202
rect 1490 31202 1619 31208
rect 1490 31192 1500 31202
rect 1660 31194 1706 31352
rect 342 31152 352 31162
rect 219 31146 352 31152
rect 858 31152 868 31162
rect 1660 31160 1666 31194
rect 1700 31160 1706 31194
rect 858 31146 1619 31152
rect 219 31112 231 31146
rect 1607 31112 1619 31146
rect 219 31106 352 31112
rect 132 31064 138 31098
rect 172 31064 178 31098
rect 342 31096 352 31106
rect 858 31106 1619 31112
rect 858 31096 868 31106
rect 132 30906 178 31064
rect 970 31056 980 31066
rect 219 31050 980 31056
rect 1490 31056 1500 31066
rect 1490 31050 1619 31056
rect 219 31016 231 31050
rect 1607 31016 1619 31050
rect 219 31010 980 31016
rect 970 31000 980 31010
rect 1490 31010 1619 31016
rect 1490 31000 1500 31010
rect 1660 31002 1706 31160
rect 342 30960 352 30970
rect 219 30954 352 30960
rect 858 30960 868 30970
rect 1660 30968 1666 31002
rect 1700 30968 1706 31002
rect 858 30954 1619 30960
rect 219 30920 231 30954
rect 1607 30920 1619 30954
rect 219 30914 352 30920
rect 132 30872 138 30906
rect 172 30872 178 30906
rect 342 30904 352 30914
rect 858 30914 1619 30920
rect 858 30904 868 30914
rect 132 30714 178 30872
rect 970 30864 980 30874
rect 219 30858 980 30864
rect 1490 30864 1500 30874
rect 1490 30858 1619 30864
rect 219 30824 231 30858
rect 1607 30824 1619 30858
rect 219 30818 980 30824
rect 970 30808 980 30818
rect 1490 30818 1619 30824
rect 1490 30808 1500 30818
rect 1660 30810 1706 30968
rect 342 30768 352 30778
rect 219 30762 352 30768
rect 858 30768 868 30778
rect 1660 30776 1666 30810
rect 1700 30776 1706 30810
rect 858 30762 1619 30768
rect 219 30728 231 30762
rect 1607 30728 1619 30762
rect 219 30722 352 30728
rect 132 30680 138 30714
rect 172 30680 178 30714
rect 342 30712 352 30722
rect 858 30722 1619 30728
rect 858 30712 868 30722
rect 132 30522 178 30680
rect 970 30672 980 30682
rect 219 30666 980 30672
rect 1490 30672 1500 30682
rect 1490 30666 1619 30672
rect 219 30632 231 30666
rect 1607 30632 1619 30666
rect 219 30626 980 30632
rect 970 30616 980 30626
rect 1490 30626 1619 30632
rect 1490 30616 1500 30626
rect 1660 30618 1706 30776
rect 342 30576 352 30586
rect 219 30570 352 30576
rect 858 30576 868 30586
rect 1660 30584 1666 30618
rect 1700 30584 1706 30618
rect 858 30570 1619 30576
rect 219 30536 231 30570
rect 1607 30536 1619 30570
rect 219 30530 352 30536
rect 132 30488 138 30522
rect 172 30488 178 30522
rect 342 30520 352 30530
rect 858 30530 1619 30536
rect 858 30520 868 30530
rect 132 30330 178 30488
rect 970 30480 980 30490
rect 219 30474 980 30480
rect 1490 30480 1500 30490
rect 1490 30474 1619 30480
rect 219 30440 231 30474
rect 1607 30440 1619 30474
rect 219 30434 980 30440
rect 970 30424 980 30434
rect 1490 30434 1619 30440
rect 1490 30424 1500 30434
rect 1660 30426 1706 30584
rect 342 30384 352 30394
rect 219 30378 352 30384
rect 858 30384 868 30394
rect 1660 30392 1666 30426
rect 1700 30392 1706 30426
rect 858 30378 1619 30384
rect 219 30344 231 30378
rect 1607 30344 1619 30378
rect 219 30338 352 30344
rect 132 30296 138 30330
rect 172 30296 178 30330
rect 342 30328 352 30338
rect 858 30338 1619 30344
rect 858 30328 868 30338
rect 132 30138 178 30296
rect 970 30288 980 30298
rect 219 30282 980 30288
rect 1490 30288 1500 30298
rect 1490 30282 1619 30288
rect 219 30248 231 30282
rect 1607 30248 1619 30282
rect 219 30242 980 30248
rect 970 30232 980 30242
rect 1490 30242 1619 30248
rect 1490 30232 1500 30242
rect 1660 30234 1706 30392
rect 342 30192 352 30202
rect 219 30186 352 30192
rect 858 30192 868 30202
rect 1660 30200 1666 30234
rect 1700 30200 1706 30234
rect 858 30186 1619 30192
rect 219 30152 231 30186
rect 1607 30152 1619 30186
rect 219 30146 352 30152
rect 132 30104 138 30138
rect 172 30104 178 30138
rect 342 30136 352 30146
rect 858 30146 1619 30152
rect 858 30136 868 30146
rect 132 29946 178 30104
rect 970 30096 980 30106
rect 219 30090 980 30096
rect 1490 30096 1500 30106
rect 1490 30090 1619 30096
rect 219 30056 231 30090
rect 1607 30056 1619 30090
rect 219 30050 980 30056
rect 970 30040 980 30050
rect 1490 30050 1619 30056
rect 1490 30040 1500 30050
rect 1660 30042 1706 30200
rect 342 30000 352 30010
rect 219 29994 352 30000
rect 858 30000 868 30010
rect 1660 30008 1666 30042
rect 1700 30008 1706 30042
rect 858 29994 1619 30000
rect 219 29960 231 29994
rect 1607 29960 1619 29994
rect 219 29954 352 29960
rect 132 29912 138 29946
rect 172 29912 178 29946
rect 342 29944 352 29954
rect 858 29954 1619 29960
rect 858 29944 868 29954
rect 132 29754 178 29912
rect 970 29904 980 29914
rect 219 29898 980 29904
rect 1490 29904 1500 29914
rect 1490 29898 1619 29904
rect 219 29864 231 29898
rect 1607 29864 1619 29898
rect 219 29858 980 29864
rect 970 29848 980 29858
rect 1490 29858 1619 29864
rect 1490 29848 1500 29858
rect 1660 29850 1706 30008
rect 342 29808 352 29818
rect 219 29802 352 29808
rect 858 29808 868 29818
rect 1660 29816 1666 29850
rect 1700 29816 1706 29850
rect 858 29802 1619 29808
rect 219 29768 231 29802
rect 1607 29768 1619 29802
rect 219 29762 352 29768
rect 132 29720 138 29754
rect 172 29720 178 29754
rect 342 29752 352 29762
rect 858 29762 1619 29768
rect 858 29752 868 29762
rect 132 29562 178 29720
rect 970 29712 980 29722
rect 219 29706 980 29712
rect 1490 29712 1500 29722
rect 1490 29706 1619 29712
rect 219 29672 231 29706
rect 1607 29672 1619 29706
rect 219 29666 980 29672
rect 970 29656 980 29666
rect 1490 29666 1619 29672
rect 1490 29656 1500 29666
rect 1660 29658 1706 29816
rect 342 29616 352 29626
rect 219 29610 352 29616
rect 858 29616 868 29626
rect 1660 29624 1666 29658
rect 1700 29624 1706 29658
rect 858 29610 1619 29616
rect 219 29576 231 29610
rect 1607 29576 1619 29610
rect 219 29570 352 29576
rect 132 29528 138 29562
rect 172 29528 178 29562
rect 342 29560 352 29570
rect 858 29570 1619 29576
rect 858 29560 868 29570
rect 132 29370 178 29528
rect 970 29520 980 29530
rect 219 29514 980 29520
rect 1490 29520 1500 29530
rect 1490 29514 1619 29520
rect 219 29480 231 29514
rect 1607 29480 1619 29514
rect 219 29474 980 29480
rect 970 29464 980 29474
rect 1490 29474 1619 29480
rect 1490 29464 1500 29474
rect 1660 29466 1706 29624
rect 342 29424 352 29434
rect 219 29418 352 29424
rect 858 29424 868 29434
rect 1660 29432 1666 29466
rect 1700 29432 1706 29466
rect 858 29418 1619 29424
rect 219 29384 231 29418
rect 1607 29384 1619 29418
rect 219 29378 352 29384
rect 132 29336 138 29370
rect 172 29336 178 29370
rect 342 29368 352 29378
rect 858 29378 1619 29384
rect 858 29368 868 29378
rect 132 29178 178 29336
rect 970 29328 980 29338
rect 219 29322 980 29328
rect 1490 29328 1500 29338
rect 1490 29322 1619 29328
rect 219 29288 231 29322
rect 1607 29288 1619 29322
rect 219 29282 980 29288
rect 970 29272 980 29282
rect 1490 29282 1619 29288
rect 1490 29272 1500 29282
rect 1660 29274 1706 29432
rect 342 29232 352 29242
rect 219 29226 352 29232
rect 858 29232 868 29242
rect 1660 29240 1666 29274
rect 1700 29240 1706 29274
rect 858 29226 1619 29232
rect 219 29192 231 29226
rect 1607 29192 1619 29226
rect 219 29186 352 29192
rect 132 29144 138 29178
rect 172 29144 178 29178
rect 342 29176 352 29186
rect 858 29186 1619 29192
rect 858 29176 868 29186
rect 132 28986 178 29144
rect 970 29136 980 29146
rect 219 29130 980 29136
rect 1490 29136 1500 29146
rect 1490 29130 1619 29136
rect 219 29096 231 29130
rect 1607 29096 1619 29130
rect 219 29090 980 29096
rect 970 29080 980 29090
rect 1490 29090 1619 29096
rect 1490 29080 1500 29090
rect 1660 29082 1706 29240
rect 342 29040 352 29050
rect 219 29034 352 29040
rect 858 29040 868 29050
rect 1660 29048 1666 29082
rect 1700 29048 1706 29082
rect 858 29034 1619 29040
rect 219 29000 231 29034
rect 1607 29000 1619 29034
rect 219 28994 352 29000
rect 132 28952 138 28986
rect 172 28952 178 28986
rect 342 28984 352 28994
rect 858 28994 1619 29000
rect 858 28984 868 28994
rect 132 28794 178 28952
rect 970 28944 980 28954
rect 219 28938 980 28944
rect 1490 28944 1500 28954
rect 1490 28938 1619 28944
rect 219 28904 231 28938
rect 1607 28904 1619 28938
rect 219 28898 980 28904
rect 970 28888 980 28898
rect 1490 28898 1619 28904
rect 1490 28888 1500 28898
rect 1660 28890 1706 29048
rect 342 28848 352 28858
rect 219 28842 352 28848
rect 858 28848 868 28858
rect 1660 28856 1666 28890
rect 1700 28856 1706 28890
rect 858 28842 1619 28848
rect 219 28808 231 28842
rect 1607 28808 1619 28842
rect 219 28802 352 28808
rect 132 28760 138 28794
rect 172 28760 178 28794
rect 342 28792 352 28802
rect 858 28802 1619 28808
rect 858 28792 868 28802
rect 132 28602 178 28760
rect 970 28752 980 28762
rect 219 28746 980 28752
rect 1490 28752 1500 28762
rect 1490 28746 1619 28752
rect 219 28712 231 28746
rect 1607 28712 1619 28746
rect 219 28706 980 28712
rect 970 28696 980 28706
rect 1490 28706 1619 28712
rect 1490 28696 1500 28706
rect 1660 28698 1706 28856
rect 342 28656 352 28666
rect 219 28650 352 28656
rect 858 28656 868 28666
rect 1660 28664 1666 28698
rect 1700 28664 1706 28698
rect 858 28650 1619 28656
rect 219 28616 231 28650
rect 1607 28616 1619 28650
rect 219 28610 352 28616
rect 132 28568 138 28602
rect 172 28568 178 28602
rect 342 28600 352 28610
rect 858 28610 1619 28616
rect 858 28600 868 28610
rect 132 28410 178 28568
rect 970 28560 980 28570
rect 219 28554 980 28560
rect 1490 28560 1500 28570
rect 1490 28554 1619 28560
rect 219 28520 231 28554
rect 1607 28520 1619 28554
rect 219 28514 980 28520
rect 970 28504 980 28514
rect 1490 28514 1619 28520
rect 1490 28504 1500 28514
rect 1660 28506 1706 28664
rect 342 28464 352 28474
rect 219 28458 352 28464
rect 858 28464 868 28474
rect 1660 28472 1666 28506
rect 1700 28472 1706 28506
rect 858 28458 1619 28464
rect 219 28424 231 28458
rect 1607 28424 1619 28458
rect 219 28418 352 28424
rect 132 28376 138 28410
rect 172 28376 178 28410
rect 342 28408 352 28418
rect 858 28418 1619 28424
rect 858 28408 868 28418
rect 132 28218 178 28376
rect 970 28368 980 28378
rect 219 28362 980 28368
rect 1490 28368 1500 28378
rect 1490 28362 1619 28368
rect 219 28328 231 28362
rect 1607 28328 1619 28362
rect 219 28322 980 28328
rect 970 28312 980 28322
rect 1490 28322 1619 28328
rect 1490 28312 1500 28322
rect 1660 28314 1706 28472
rect 342 28272 352 28282
rect 219 28266 352 28272
rect 858 28272 868 28282
rect 1660 28280 1666 28314
rect 1700 28280 1706 28314
rect 858 28266 1619 28272
rect 219 28232 231 28266
rect 1607 28232 1619 28266
rect 219 28226 352 28232
rect 132 28184 138 28218
rect 172 28184 178 28218
rect 342 28216 352 28226
rect 858 28226 1619 28232
rect 858 28216 868 28226
rect 132 28026 178 28184
rect 970 28176 980 28186
rect 219 28170 980 28176
rect 1490 28176 1500 28186
rect 1490 28170 1619 28176
rect 219 28136 231 28170
rect 1607 28136 1619 28170
rect 219 28130 980 28136
rect 970 28120 980 28130
rect 1490 28130 1619 28136
rect 1490 28120 1500 28130
rect 1660 28122 1706 28280
rect 342 28080 352 28090
rect 219 28074 352 28080
rect 858 28080 868 28090
rect 1660 28088 1666 28122
rect 1700 28088 1706 28122
rect 858 28074 1619 28080
rect 219 28040 231 28074
rect 1607 28040 1619 28074
rect 219 28034 352 28040
rect 132 27992 138 28026
rect 172 27992 178 28026
rect 342 28024 352 28034
rect 858 28034 1619 28040
rect 858 28024 868 28034
rect 132 27834 178 27992
rect 970 27984 980 27994
rect 219 27978 980 27984
rect 1490 27984 1500 27994
rect 1490 27978 1619 27984
rect 219 27944 231 27978
rect 1607 27944 1619 27978
rect 219 27938 980 27944
rect 970 27928 980 27938
rect 1490 27938 1619 27944
rect 1490 27928 1500 27938
rect 1660 27930 1706 28088
rect 342 27888 352 27898
rect 219 27882 352 27888
rect 858 27888 868 27898
rect 1660 27896 1666 27930
rect 1700 27896 1706 27930
rect 858 27882 1619 27888
rect 219 27848 231 27882
rect 1607 27848 1619 27882
rect 219 27842 352 27848
rect 132 27800 138 27834
rect 172 27800 178 27834
rect 342 27832 352 27842
rect 858 27842 1619 27848
rect 858 27832 868 27842
rect 132 27642 178 27800
rect 970 27792 980 27802
rect 219 27786 980 27792
rect 1490 27792 1500 27802
rect 1490 27786 1619 27792
rect 219 27752 231 27786
rect 1607 27752 1619 27786
rect 219 27746 980 27752
rect 970 27736 980 27746
rect 1490 27746 1619 27752
rect 1490 27736 1500 27746
rect 1660 27738 1706 27896
rect 342 27696 352 27706
rect 219 27690 352 27696
rect 858 27696 868 27706
rect 1660 27704 1666 27738
rect 1700 27704 1706 27738
rect 858 27690 1619 27696
rect 219 27656 231 27690
rect 1607 27656 1619 27690
rect 219 27650 352 27656
rect 132 27608 138 27642
rect 172 27608 178 27642
rect 342 27640 352 27650
rect 858 27650 1619 27656
rect 858 27640 868 27650
rect 132 27450 178 27608
rect 970 27600 980 27610
rect 219 27594 980 27600
rect 1490 27600 1500 27610
rect 1490 27594 1619 27600
rect 219 27560 231 27594
rect 1607 27560 1619 27594
rect 219 27554 980 27560
rect 970 27544 980 27554
rect 1490 27554 1619 27560
rect 1490 27544 1500 27554
rect 1660 27546 1706 27704
rect 342 27504 352 27514
rect 219 27498 352 27504
rect 858 27504 868 27514
rect 1660 27512 1666 27546
rect 1700 27512 1706 27546
rect 858 27498 1619 27504
rect 219 27464 231 27498
rect 1607 27464 1619 27498
rect 219 27458 352 27464
rect 132 27416 138 27450
rect 172 27416 178 27450
rect 342 27448 352 27458
rect 858 27458 1619 27464
rect 858 27448 868 27458
rect 132 27258 178 27416
rect 970 27408 980 27418
rect 219 27402 980 27408
rect 1490 27408 1500 27418
rect 1490 27402 1619 27408
rect 219 27368 231 27402
rect 1607 27368 1619 27402
rect 219 27362 980 27368
rect 970 27352 980 27362
rect 1490 27362 1619 27368
rect 1490 27352 1500 27362
rect 1660 27354 1706 27512
rect 342 27312 352 27322
rect 219 27306 352 27312
rect 858 27312 868 27322
rect 1660 27320 1666 27354
rect 1700 27320 1706 27354
rect 858 27306 1619 27312
rect 219 27272 231 27306
rect 1607 27272 1619 27306
rect 219 27266 352 27272
rect 132 27224 138 27258
rect 172 27224 178 27258
rect 342 27256 352 27266
rect 858 27266 1619 27272
rect 858 27256 868 27266
rect 132 27066 178 27224
rect 970 27216 980 27226
rect 219 27210 980 27216
rect 1490 27216 1500 27226
rect 1490 27210 1619 27216
rect 219 27176 231 27210
rect 1607 27176 1619 27210
rect 219 27170 980 27176
rect 970 27160 980 27170
rect 1490 27170 1619 27176
rect 1490 27160 1500 27170
rect 1660 27162 1706 27320
rect 342 27120 352 27130
rect 219 27114 352 27120
rect 858 27120 868 27130
rect 1660 27128 1666 27162
rect 1700 27128 1706 27162
rect 858 27114 1619 27120
rect 219 27080 231 27114
rect 1607 27080 1619 27114
rect 219 27074 352 27080
rect 132 27032 138 27066
rect 172 27032 178 27066
rect 342 27064 352 27074
rect 858 27074 1619 27080
rect 858 27064 868 27074
rect 132 26874 178 27032
rect 970 27024 980 27034
rect 219 27018 980 27024
rect 1490 27024 1500 27034
rect 1490 27018 1619 27024
rect 219 26984 231 27018
rect 1607 26984 1619 27018
rect 219 26978 980 26984
rect 970 26968 980 26978
rect 1490 26978 1619 26984
rect 1490 26968 1500 26978
rect 1660 26970 1706 27128
rect 342 26928 352 26938
rect 219 26922 352 26928
rect 858 26928 868 26938
rect 1660 26936 1666 26970
rect 1700 26936 1706 26970
rect 858 26922 1619 26928
rect 219 26888 231 26922
rect 1607 26888 1619 26922
rect 219 26882 352 26888
rect 132 26840 138 26874
rect 172 26840 178 26874
rect 342 26872 352 26882
rect 858 26882 1619 26888
rect 858 26872 868 26882
rect 132 26682 178 26840
rect 970 26832 980 26842
rect 219 26826 980 26832
rect 1490 26832 1500 26842
rect 1490 26826 1619 26832
rect 219 26792 231 26826
rect 1607 26792 1619 26826
rect 219 26786 980 26792
rect 970 26776 980 26786
rect 1490 26786 1619 26792
rect 1490 26776 1500 26786
rect 1660 26778 1706 26936
rect 342 26736 352 26746
rect 219 26730 352 26736
rect 858 26736 868 26746
rect 1660 26744 1666 26778
rect 1700 26744 1706 26778
rect 858 26730 1619 26736
rect 219 26696 231 26730
rect 1607 26696 1619 26730
rect 219 26690 352 26696
rect 132 26648 138 26682
rect 172 26648 178 26682
rect 342 26680 352 26690
rect 858 26690 1619 26696
rect 858 26680 868 26690
rect 132 26490 178 26648
rect 970 26640 980 26650
rect 219 26634 980 26640
rect 1490 26640 1500 26650
rect 1490 26634 1619 26640
rect 219 26600 231 26634
rect 1607 26600 1619 26634
rect 219 26594 980 26600
rect 970 26584 980 26594
rect 1490 26594 1619 26600
rect 1490 26584 1500 26594
rect 1660 26586 1706 26744
rect 342 26544 352 26554
rect 219 26538 352 26544
rect 858 26544 868 26554
rect 1660 26552 1666 26586
rect 1700 26552 1706 26586
rect 858 26538 1619 26544
rect 219 26504 231 26538
rect 1607 26504 1619 26538
rect 219 26498 352 26504
rect 132 26456 138 26490
rect 172 26456 178 26490
rect 342 26488 352 26498
rect 858 26498 1619 26504
rect 858 26488 868 26498
rect 132 26298 178 26456
rect 970 26448 980 26458
rect 219 26442 980 26448
rect 1490 26448 1500 26458
rect 1490 26442 1619 26448
rect 219 26408 231 26442
rect 1607 26408 1619 26442
rect 219 26402 980 26408
rect 970 26392 980 26402
rect 1490 26402 1619 26408
rect 1490 26392 1500 26402
rect 1660 26394 1706 26552
rect 342 26352 352 26362
rect 219 26346 352 26352
rect 858 26352 868 26362
rect 1660 26360 1666 26394
rect 1700 26360 1706 26394
rect 858 26346 1619 26352
rect 219 26312 231 26346
rect 1607 26312 1619 26346
rect 219 26306 352 26312
rect 132 26264 138 26298
rect 172 26264 178 26298
rect 342 26296 352 26306
rect 858 26306 1619 26312
rect 858 26296 868 26306
rect 132 26106 178 26264
rect 970 26256 980 26266
rect 219 26250 980 26256
rect 1490 26256 1500 26266
rect 1490 26250 1619 26256
rect 219 26216 231 26250
rect 1607 26216 1619 26250
rect 219 26210 980 26216
rect 970 26200 980 26210
rect 1490 26210 1619 26216
rect 1490 26200 1500 26210
rect 1660 26202 1706 26360
rect 342 26160 352 26170
rect 219 26154 352 26160
rect 858 26160 868 26170
rect 1660 26168 1666 26202
rect 1700 26168 1706 26202
rect 858 26154 1619 26160
rect 219 26120 231 26154
rect 1607 26120 1619 26154
rect 219 26114 352 26120
rect 132 26072 138 26106
rect 172 26072 178 26106
rect 342 26104 352 26114
rect 858 26114 1619 26120
rect 858 26104 868 26114
rect 132 25914 178 26072
rect 970 26064 980 26074
rect 219 26058 980 26064
rect 1490 26064 1500 26074
rect 1490 26058 1619 26064
rect 219 26024 231 26058
rect 1607 26024 1619 26058
rect 219 26018 980 26024
rect 970 26008 980 26018
rect 1490 26018 1619 26024
rect 1490 26008 1500 26018
rect 1660 26010 1706 26168
rect 342 25968 352 25978
rect 219 25962 352 25968
rect 858 25968 868 25978
rect 1660 25976 1666 26010
rect 1700 25976 1706 26010
rect 858 25962 1619 25968
rect 219 25928 231 25962
rect 1607 25928 1619 25962
rect 219 25922 352 25928
rect 132 25880 138 25914
rect 172 25880 178 25914
rect 342 25912 352 25922
rect 858 25922 1619 25928
rect 858 25912 868 25922
rect 132 25722 178 25880
rect 970 25872 980 25882
rect 219 25866 980 25872
rect 1490 25872 1500 25882
rect 1490 25866 1619 25872
rect 219 25832 231 25866
rect 1607 25832 1619 25866
rect 219 25826 980 25832
rect 970 25816 980 25826
rect 1490 25826 1619 25832
rect 1490 25816 1500 25826
rect 1660 25818 1706 25976
rect 342 25776 352 25786
rect 219 25770 352 25776
rect 858 25776 868 25786
rect 1660 25784 1666 25818
rect 1700 25784 1706 25818
rect 858 25770 1619 25776
rect 219 25736 231 25770
rect 1607 25736 1619 25770
rect 219 25730 352 25736
rect 132 25688 138 25722
rect 172 25688 178 25722
rect 342 25720 352 25730
rect 858 25730 1619 25736
rect 858 25720 868 25730
rect 132 25530 178 25688
rect 970 25680 980 25690
rect 219 25674 980 25680
rect 1490 25680 1500 25690
rect 1490 25674 1619 25680
rect 219 25640 231 25674
rect 1607 25640 1619 25674
rect 219 25634 980 25640
rect 970 25624 980 25634
rect 1490 25634 1619 25640
rect 1490 25624 1500 25634
rect 1660 25626 1706 25784
rect 342 25584 352 25594
rect 219 25578 352 25584
rect 858 25584 868 25594
rect 1660 25592 1666 25626
rect 1700 25592 1706 25626
rect 858 25578 1619 25584
rect 219 25544 231 25578
rect 1607 25544 1619 25578
rect 219 25538 352 25544
rect 132 25496 138 25530
rect 172 25496 178 25530
rect 342 25528 352 25538
rect 858 25538 1619 25544
rect 858 25528 868 25538
rect 132 25338 178 25496
rect 970 25488 980 25498
rect 219 25482 980 25488
rect 1490 25488 1500 25498
rect 1490 25482 1619 25488
rect 219 25448 231 25482
rect 1607 25448 1619 25482
rect 219 25442 980 25448
rect 970 25432 980 25442
rect 1490 25442 1619 25448
rect 1490 25432 1500 25442
rect 1660 25434 1706 25592
rect 342 25392 352 25402
rect 219 25386 352 25392
rect 858 25392 868 25402
rect 1660 25400 1666 25434
rect 1700 25400 1706 25434
rect 858 25386 1619 25392
rect 219 25352 231 25386
rect 1607 25352 1619 25386
rect 219 25346 352 25352
rect 132 25304 138 25338
rect 172 25304 178 25338
rect 342 25336 352 25346
rect 858 25346 1619 25352
rect 858 25336 868 25346
rect 132 25146 178 25304
rect 970 25296 980 25306
rect 219 25290 980 25296
rect 1490 25296 1500 25306
rect 1490 25290 1619 25296
rect 219 25256 231 25290
rect 1607 25256 1619 25290
rect 219 25250 980 25256
rect 970 25240 980 25250
rect 1490 25250 1619 25256
rect 1490 25240 1500 25250
rect 1660 25242 1706 25400
rect 342 25200 352 25210
rect 219 25194 352 25200
rect 858 25200 868 25210
rect 1660 25208 1666 25242
rect 1700 25208 1706 25242
rect 858 25194 1619 25200
rect 219 25160 231 25194
rect 1607 25160 1619 25194
rect 219 25154 352 25160
rect 132 25112 138 25146
rect 172 25112 178 25146
rect 342 25144 352 25154
rect 858 25154 1619 25160
rect 858 25144 868 25154
rect 132 24954 178 25112
rect 970 25104 980 25114
rect 219 25098 980 25104
rect 1490 25104 1500 25114
rect 1490 25098 1619 25104
rect 219 25064 231 25098
rect 1607 25064 1619 25098
rect 219 25058 980 25064
rect 970 25048 980 25058
rect 1490 25058 1619 25064
rect 1490 25048 1500 25058
rect 1660 25050 1706 25208
rect 342 25008 352 25018
rect 219 25002 352 25008
rect 858 25008 868 25018
rect 1660 25016 1666 25050
rect 1700 25016 1706 25050
rect 858 25002 1619 25008
rect 219 24968 231 25002
rect 1607 24968 1619 25002
rect 219 24962 352 24968
rect 132 24920 138 24954
rect 172 24920 178 24954
rect 342 24952 352 24962
rect 858 24962 1619 24968
rect 858 24952 868 24962
rect 132 24762 178 24920
rect 970 24912 980 24922
rect 219 24906 980 24912
rect 1490 24912 1500 24922
rect 1490 24906 1619 24912
rect 219 24872 231 24906
rect 1607 24872 1619 24906
rect 219 24866 980 24872
rect 970 24856 980 24866
rect 1490 24866 1619 24872
rect 1490 24856 1500 24866
rect 1660 24858 1706 25016
rect 342 24816 352 24826
rect 219 24810 352 24816
rect 858 24816 868 24826
rect 1660 24824 1666 24858
rect 1700 24824 1706 24858
rect 858 24810 1619 24816
rect 219 24776 231 24810
rect 1607 24776 1619 24810
rect 219 24770 352 24776
rect 132 24728 138 24762
rect 172 24728 178 24762
rect 342 24760 352 24770
rect 858 24770 1619 24776
rect 858 24760 868 24770
rect 132 24570 178 24728
rect 970 24720 980 24730
rect 219 24714 980 24720
rect 1490 24720 1500 24730
rect 1490 24714 1619 24720
rect 219 24680 231 24714
rect 1607 24680 1619 24714
rect 219 24674 980 24680
rect 970 24664 980 24674
rect 1490 24674 1619 24680
rect 1490 24664 1500 24674
rect 1660 24666 1706 24824
rect 342 24624 352 24634
rect 219 24618 352 24624
rect 858 24624 868 24634
rect 1660 24632 1666 24666
rect 1700 24632 1706 24666
rect 858 24618 1619 24624
rect 219 24584 231 24618
rect 1607 24584 1619 24618
rect 219 24578 352 24584
rect 132 24536 138 24570
rect 172 24536 178 24570
rect 342 24568 352 24578
rect 858 24578 1619 24584
rect 858 24568 868 24578
rect 132 24378 178 24536
rect 970 24528 980 24538
rect 219 24522 980 24528
rect 1490 24528 1500 24538
rect 1490 24522 1619 24528
rect 219 24488 231 24522
rect 1607 24488 1619 24522
rect 219 24482 980 24488
rect 970 24472 980 24482
rect 1490 24482 1619 24488
rect 1490 24472 1500 24482
rect 1660 24474 1706 24632
rect 342 24432 352 24442
rect 219 24426 352 24432
rect 858 24432 868 24442
rect 1660 24440 1666 24474
rect 1700 24440 1706 24474
rect 858 24426 1619 24432
rect 219 24392 231 24426
rect 1607 24392 1619 24426
rect 219 24386 352 24392
rect 132 24344 138 24378
rect 172 24344 178 24378
rect 342 24376 352 24386
rect 858 24386 1619 24392
rect 858 24376 868 24386
rect 132 24186 178 24344
rect 970 24336 980 24346
rect 219 24330 980 24336
rect 1490 24336 1500 24346
rect 1490 24330 1619 24336
rect 219 24296 231 24330
rect 1607 24296 1619 24330
rect 219 24290 980 24296
rect 970 24280 980 24290
rect 1490 24290 1619 24296
rect 1490 24280 1500 24290
rect 1660 24282 1706 24440
rect 342 24240 352 24250
rect 219 24234 352 24240
rect 858 24240 868 24250
rect 1660 24248 1666 24282
rect 1700 24248 1706 24282
rect 858 24234 1619 24240
rect 219 24200 231 24234
rect 1607 24200 1619 24234
rect 219 24194 352 24200
rect 132 24152 138 24186
rect 172 24152 178 24186
rect 342 24184 352 24194
rect 858 24194 1619 24200
rect 858 24184 868 24194
rect 132 23994 178 24152
rect 970 24144 980 24154
rect 219 24138 980 24144
rect 1490 24144 1500 24154
rect 1490 24138 1619 24144
rect 219 24104 231 24138
rect 1607 24104 1619 24138
rect 219 24098 980 24104
rect 970 24088 980 24098
rect 1490 24098 1619 24104
rect 1490 24088 1500 24098
rect 1660 24090 1706 24248
rect 342 24048 352 24058
rect 219 24042 352 24048
rect 858 24048 868 24058
rect 1660 24056 1666 24090
rect 1700 24056 1706 24090
rect 858 24042 1619 24048
rect 219 24008 231 24042
rect 1607 24008 1619 24042
rect 219 24002 352 24008
rect 132 23960 138 23994
rect 172 23960 178 23994
rect 342 23992 352 24002
rect 858 24002 1619 24008
rect 858 23992 868 24002
rect 132 23802 178 23960
rect 970 23952 980 23962
rect 219 23946 980 23952
rect 1490 23952 1500 23962
rect 1490 23946 1619 23952
rect 219 23912 231 23946
rect 1607 23912 1619 23946
rect 219 23906 980 23912
rect 970 23896 980 23906
rect 1490 23906 1619 23912
rect 1490 23896 1500 23906
rect 1660 23898 1706 24056
rect 342 23856 352 23866
rect 219 23850 352 23856
rect 858 23856 868 23866
rect 1660 23864 1666 23898
rect 1700 23864 1706 23898
rect 858 23850 1619 23856
rect 219 23816 231 23850
rect 1607 23816 1619 23850
rect 219 23810 352 23816
rect 132 23768 138 23802
rect 172 23768 178 23802
rect 342 23800 352 23810
rect 858 23810 1619 23816
rect 858 23800 868 23810
rect 132 23610 178 23768
rect 970 23760 980 23770
rect 219 23754 980 23760
rect 1490 23760 1500 23770
rect 1490 23754 1619 23760
rect 219 23720 231 23754
rect 1607 23720 1619 23754
rect 219 23714 980 23720
rect 970 23704 980 23714
rect 1490 23714 1619 23720
rect 1490 23704 1500 23714
rect 1660 23706 1706 23864
rect 342 23664 352 23674
rect 219 23658 352 23664
rect 858 23664 868 23674
rect 1660 23672 1666 23706
rect 1700 23672 1706 23706
rect 858 23658 1619 23664
rect 219 23624 231 23658
rect 1607 23624 1619 23658
rect 219 23618 352 23624
rect 132 23576 138 23610
rect 172 23576 178 23610
rect 342 23608 352 23618
rect 858 23618 1619 23624
rect 858 23608 868 23618
rect 132 23418 178 23576
rect 970 23568 980 23578
rect 219 23562 980 23568
rect 1490 23568 1500 23578
rect 1490 23562 1619 23568
rect 219 23528 231 23562
rect 1607 23528 1619 23562
rect 219 23522 980 23528
rect 970 23512 980 23522
rect 1490 23522 1619 23528
rect 1490 23512 1500 23522
rect 1660 23514 1706 23672
rect 342 23472 352 23482
rect 219 23466 352 23472
rect 858 23472 868 23482
rect 1660 23480 1666 23514
rect 1700 23480 1706 23514
rect 858 23466 1619 23472
rect 219 23432 231 23466
rect 1607 23432 1619 23466
rect 219 23426 352 23432
rect 132 23384 138 23418
rect 172 23384 178 23418
rect 342 23416 352 23426
rect 858 23426 1619 23432
rect 858 23416 868 23426
rect 132 23226 178 23384
rect 970 23376 980 23386
rect 219 23370 980 23376
rect 1490 23376 1500 23386
rect 1490 23370 1619 23376
rect 219 23336 231 23370
rect 1607 23336 1619 23370
rect 219 23330 980 23336
rect 970 23320 980 23330
rect 1490 23330 1619 23336
rect 1490 23320 1500 23330
rect 1660 23322 1706 23480
rect 342 23280 352 23290
rect 219 23274 352 23280
rect 858 23280 868 23290
rect 1660 23288 1666 23322
rect 1700 23288 1706 23322
rect 858 23274 1619 23280
rect 219 23240 231 23274
rect 1607 23240 1619 23274
rect 219 23234 352 23240
rect 132 23192 138 23226
rect 172 23192 178 23226
rect 342 23224 352 23234
rect 858 23234 1619 23240
rect 858 23224 868 23234
rect 132 21656 178 23192
rect 970 23184 980 23194
rect 219 23178 980 23184
rect 1490 23184 1500 23194
rect 1490 23178 1619 23184
rect 219 23144 231 23178
rect 1607 23144 1619 23178
rect 219 23138 980 23144
rect 970 23128 980 23138
rect 1490 23138 1619 23144
rect 1660 23168 1706 23288
rect 1490 23128 1500 23138
rect 1660 23130 1708 23168
rect 342 23088 352 23098
rect 219 23082 352 23088
rect 858 23088 868 23098
rect 1660 23096 1666 23130
rect 1700 23096 1708 23130
rect 858 23082 1619 23088
rect 219 23048 231 23082
rect 1607 23048 1619 23082
rect 219 23042 352 23048
rect 342 23032 352 23042
rect 858 23042 1619 23048
rect 858 23032 868 23042
rect 334 22768 876 22780
rect 330 21986 340 22768
rect 870 21986 880 22768
rect 334 21974 876 21986
rect 342 21710 352 21720
rect 219 21704 352 21710
rect 858 21710 868 21720
rect 858 21704 1619 21710
rect 219 21670 231 21704
rect 1607 21670 1619 21704
rect 219 21664 352 21670
rect 132 21622 138 21656
rect 172 21622 178 21656
rect 342 21654 352 21664
rect 858 21664 1619 21670
rect 858 21654 868 21664
rect 132 21464 178 21622
rect 970 21614 980 21624
rect 219 21608 980 21614
rect 1490 21614 1500 21624
rect 1490 21608 1619 21614
rect 219 21574 231 21608
rect 1607 21574 1619 21608
rect 219 21568 980 21574
rect 970 21558 980 21568
rect 1490 21568 1619 21574
rect 1490 21558 1500 21568
rect 1660 21560 1708 23096
rect 342 21518 352 21528
rect 219 21512 352 21518
rect 858 21518 868 21528
rect 1660 21526 1666 21560
rect 1700 21526 1708 21560
rect 858 21512 1619 21518
rect 219 21478 231 21512
rect 1607 21478 1619 21512
rect 219 21472 352 21478
rect 132 21430 138 21464
rect 172 21430 178 21464
rect 342 21462 352 21472
rect 858 21472 1619 21478
rect 858 21462 868 21472
rect 132 21272 178 21430
rect 970 21422 980 21432
rect 219 21416 980 21422
rect 1490 21422 1500 21432
rect 1490 21416 1619 21422
rect 219 21382 231 21416
rect 1607 21382 1619 21416
rect 219 21376 980 21382
rect 970 21366 980 21376
rect 1490 21376 1619 21382
rect 1490 21366 1500 21376
rect 1660 21368 1708 21526
rect 342 21326 352 21336
rect 219 21320 352 21326
rect 858 21326 868 21336
rect 1660 21334 1666 21368
rect 1700 21334 1708 21368
rect 858 21320 1619 21326
rect 219 21286 231 21320
rect 1607 21286 1619 21320
rect 219 21280 352 21286
rect 132 21238 138 21272
rect 172 21238 178 21272
rect 342 21270 352 21280
rect 858 21280 1619 21286
rect 858 21270 868 21280
rect 132 21080 178 21238
rect 970 21230 980 21240
rect 219 21224 980 21230
rect 1490 21230 1500 21240
rect 1490 21224 1619 21230
rect 219 21190 231 21224
rect 1607 21190 1619 21224
rect 219 21184 980 21190
rect 970 21174 980 21184
rect 1490 21184 1619 21190
rect 1490 21174 1500 21184
rect 1660 21176 1708 21334
rect 342 21134 352 21144
rect 219 21128 352 21134
rect 858 21134 868 21144
rect 1660 21142 1666 21176
rect 1700 21142 1708 21176
rect 858 21128 1619 21134
rect 219 21094 231 21128
rect 1607 21094 1619 21128
rect 219 21088 352 21094
rect 132 21046 138 21080
rect 172 21046 178 21080
rect 342 21078 352 21088
rect 858 21088 1619 21094
rect 858 21078 868 21088
rect 132 20888 178 21046
rect 970 21038 980 21048
rect 219 21032 980 21038
rect 1490 21038 1500 21048
rect 1490 21032 1619 21038
rect 219 20998 231 21032
rect 1607 20998 1619 21032
rect 219 20992 980 20998
rect 970 20982 980 20992
rect 1490 20992 1619 20998
rect 1490 20982 1500 20992
rect 1660 20984 1708 21142
rect 342 20942 352 20952
rect 219 20936 352 20942
rect 858 20942 868 20952
rect 1660 20950 1666 20984
rect 1700 20950 1708 20984
rect 858 20936 1619 20942
rect 219 20902 231 20936
rect 1607 20902 1619 20936
rect 219 20896 352 20902
rect 132 20854 138 20888
rect 172 20854 178 20888
rect 342 20886 352 20896
rect 858 20896 1619 20902
rect 858 20886 868 20896
rect 132 20696 178 20854
rect 970 20846 980 20856
rect 219 20840 980 20846
rect 1490 20846 1500 20856
rect 1490 20840 1619 20846
rect 219 20806 231 20840
rect 1607 20806 1619 20840
rect 219 20800 980 20806
rect 970 20790 980 20800
rect 1490 20800 1619 20806
rect 1490 20790 1500 20800
rect 1660 20792 1708 20950
rect 342 20750 352 20760
rect 219 20744 352 20750
rect 858 20750 868 20760
rect 1660 20758 1666 20792
rect 1700 20758 1708 20792
rect 858 20744 1619 20750
rect 219 20710 231 20744
rect 1607 20710 1619 20744
rect 219 20704 352 20710
rect 132 20662 138 20696
rect 172 20662 178 20696
rect 342 20694 352 20704
rect 858 20704 1619 20710
rect 858 20694 868 20704
rect 132 20504 178 20662
rect 970 20654 980 20664
rect 219 20648 980 20654
rect 1490 20654 1500 20664
rect 1490 20648 1619 20654
rect 219 20614 231 20648
rect 1607 20614 1619 20648
rect 219 20608 980 20614
rect 970 20598 980 20608
rect 1490 20608 1619 20614
rect 1490 20598 1500 20608
rect 1660 20600 1708 20758
rect 342 20558 352 20568
rect 219 20552 352 20558
rect 858 20558 868 20568
rect 1660 20566 1666 20600
rect 1700 20566 1708 20600
rect 858 20552 1619 20558
rect 219 20518 231 20552
rect 1607 20518 1619 20552
rect 219 20512 352 20518
rect 132 20470 138 20504
rect 172 20470 178 20504
rect 342 20502 352 20512
rect 858 20512 1619 20518
rect 858 20502 868 20512
rect 132 20312 178 20470
rect 970 20462 980 20472
rect 219 20456 980 20462
rect 1490 20462 1500 20472
rect 1490 20456 1619 20462
rect 219 20422 231 20456
rect 1607 20422 1619 20456
rect 219 20416 980 20422
rect 970 20406 980 20416
rect 1490 20416 1619 20422
rect 1490 20406 1500 20416
rect 1660 20408 1708 20566
rect 342 20366 352 20376
rect 219 20360 352 20366
rect 858 20366 868 20376
rect 1660 20374 1666 20408
rect 1700 20374 1708 20408
rect 858 20360 1619 20366
rect 219 20326 231 20360
rect 1607 20326 1619 20360
rect 219 20320 352 20326
rect 132 20278 138 20312
rect 172 20278 178 20312
rect 342 20310 352 20320
rect 858 20320 1619 20326
rect 858 20310 868 20320
rect 132 20120 178 20278
rect 970 20270 980 20280
rect 219 20264 980 20270
rect 1490 20270 1500 20280
rect 1490 20264 1619 20270
rect 219 20230 231 20264
rect 1607 20230 1619 20264
rect 219 20224 980 20230
rect 970 20214 980 20224
rect 1490 20224 1619 20230
rect 1490 20214 1500 20224
rect 1660 20216 1708 20374
rect 342 20174 352 20184
rect 219 20168 352 20174
rect 858 20174 868 20184
rect 1660 20182 1666 20216
rect 1700 20182 1708 20216
rect 858 20168 1619 20174
rect 219 20134 231 20168
rect 1607 20134 1619 20168
rect 219 20128 352 20134
rect 132 20086 138 20120
rect 172 20086 178 20120
rect 342 20118 352 20128
rect 858 20128 1619 20134
rect 858 20118 868 20128
rect 132 19928 178 20086
rect 970 20078 980 20088
rect 219 20072 980 20078
rect 1490 20078 1500 20088
rect 1490 20072 1619 20078
rect 219 20038 231 20072
rect 1607 20038 1619 20072
rect 219 20032 980 20038
rect 970 20022 980 20032
rect 1490 20032 1619 20038
rect 1490 20022 1500 20032
rect 1660 20024 1708 20182
rect 342 19982 352 19992
rect 219 19976 352 19982
rect 858 19982 868 19992
rect 1660 19990 1666 20024
rect 1700 19990 1708 20024
rect 858 19976 1619 19982
rect 219 19942 231 19976
rect 1607 19942 1619 19976
rect 219 19936 352 19942
rect 132 19894 138 19928
rect 172 19894 178 19928
rect 342 19926 352 19936
rect 858 19936 1619 19942
rect 858 19926 868 19936
rect 132 19736 178 19894
rect 970 19886 980 19896
rect 219 19880 980 19886
rect 1490 19886 1500 19896
rect 1490 19880 1619 19886
rect 219 19846 231 19880
rect 1607 19846 1619 19880
rect 219 19840 980 19846
rect 970 19830 980 19840
rect 1490 19840 1619 19846
rect 1490 19830 1500 19840
rect 1660 19832 1708 19990
rect 342 19790 352 19800
rect 219 19784 352 19790
rect 858 19790 868 19800
rect 1660 19798 1666 19832
rect 1700 19798 1708 19832
rect 858 19784 1619 19790
rect 219 19750 231 19784
rect 1607 19750 1619 19784
rect 219 19744 352 19750
rect 132 19702 138 19736
rect 172 19702 178 19736
rect 342 19734 352 19744
rect 858 19744 1619 19750
rect 858 19734 868 19744
rect 132 19544 178 19702
rect 970 19694 980 19704
rect 219 19688 980 19694
rect 1490 19694 1500 19704
rect 1490 19688 1619 19694
rect 219 19654 231 19688
rect 1607 19654 1619 19688
rect 219 19648 980 19654
rect 970 19638 980 19648
rect 1490 19648 1619 19654
rect 1490 19638 1500 19648
rect 1660 19640 1708 19798
rect 342 19598 352 19608
rect 219 19592 352 19598
rect 858 19598 868 19608
rect 1660 19606 1666 19640
rect 1700 19606 1708 19640
rect 858 19592 1619 19598
rect 219 19558 231 19592
rect 1607 19558 1619 19592
rect 219 19552 352 19558
rect 132 19510 138 19544
rect 172 19510 178 19544
rect 342 19542 352 19552
rect 858 19552 1619 19558
rect 858 19542 868 19552
rect 132 19352 178 19510
rect 970 19502 980 19512
rect 219 19496 980 19502
rect 1490 19502 1500 19512
rect 1490 19496 1619 19502
rect 219 19462 231 19496
rect 1607 19462 1619 19496
rect 219 19456 980 19462
rect 970 19446 980 19456
rect 1490 19456 1619 19462
rect 1490 19446 1500 19456
rect 1660 19448 1708 19606
rect 342 19406 352 19416
rect 219 19400 352 19406
rect 858 19406 868 19416
rect 1660 19414 1666 19448
rect 1700 19414 1708 19448
rect 858 19400 1619 19406
rect 219 19366 231 19400
rect 1607 19366 1619 19400
rect 219 19360 352 19366
rect 132 19318 138 19352
rect 172 19318 178 19352
rect 342 19350 352 19360
rect 858 19360 1619 19366
rect 858 19350 868 19360
rect 132 19160 178 19318
rect 970 19310 980 19320
rect 219 19304 980 19310
rect 1490 19310 1500 19320
rect 1490 19304 1619 19310
rect 219 19270 231 19304
rect 1607 19270 1619 19304
rect 219 19264 980 19270
rect 970 19254 980 19264
rect 1490 19264 1619 19270
rect 1490 19254 1500 19264
rect 1660 19256 1708 19414
rect 342 19214 352 19224
rect 219 19208 352 19214
rect 858 19214 868 19224
rect 1660 19222 1666 19256
rect 1700 19222 1708 19256
rect 858 19208 1619 19214
rect 219 19174 231 19208
rect 1607 19174 1619 19208
rect 219 19168 352 19174
rect 132 19126 138 19160
rect 172 19126 178 19160
rect 342 19158 352 19168
rect 858 19168 1619 19174
rect 858 19158 868 19168
rect 132 18968 178 19126
rect 970 19118 980 19128
rect 219 19112 980 19118
rect 1490 19118 1500 19128
rect 1490 19112 1619 19118
rect 219 19078 231 19112
rect 1607 19078 1619 19112
rect 219 19072 980 19078
rect 970 19062 980 19072
rect 1490 19072 1619 19078
rect 1490 19062 1500 19072
rect 1660 19064 1708 19222
rect 342 19022 352 19032
rect 219 19016 352 19022
rect 858 19022 868 19032
rect 1660 19030 1666 19064
rect 1700 19030 1708 19064
rect 858 19016 1619 19022
rect 219 18982 231 19016
rect 1607 18982 1619 19016
rect 219 18976 352 18982
rect 132 18934 138 18968
rect 172 18934 178 18968
rect 342 18966 352 18976
rect 858 18976 1619 18982
rect 858 18966 868 18976
rect 132 18776 178 18934
rect 970 18926 980 18936
rect 219 18920 980 18926
rect 1490 18926 1500 18936
rect 1490 18920 1619 18926
rect 219 18886 231 18920
rect 1607 18886 1619 18920
rect 219 18880 980 18886
rect 970 18870 980 18880
rect 1490 18880 1619 18886
rect 1490 18870 1500 18880
rect 1660 18872 1708 19030
rect 342 18830 352 18840
rect 219 18824 352 18830
rect 858 18830 868 18840
rect 1660 18838 1666 18872
rect 1700 18838 1708 18872
rect 858 18824 1619 18830
rect 219 18790 231 18824
rect 1607 18790 1619 18824
rect 219 18784 352 18790
rect 132 18742 138 18776
rect 172 18742 178 18776
rect 342 18774 352 18784
rect 858 18784 1619 18790
rect 858 18774 868 18784
rect 132 18584 178 18742
rect 970 18734 980 18744
rect 219 18728 980 18734
rect 1490 18734 1500 18744
rect 1490 18728 1619 18734
rect 219 18694 231 18728
rect 1607 18694 1619 18728
rect 219 18688 980 18694
rect 970 18678 980 18688
rect 1490 18688 1619 18694
rect 1490 18678 1500 18688
rect 1660 18680 1708 18838
rect 342 18638 352 18648
rect 219 18632 352 18638
rect 858 18638 868 18648
rect 1660 18646 1666 18680
rect 1700 18646 1708 18680
rect 858 18632 1619 18638
rect 219 18598 231 18632
rect 1607 18598 1619 18632
rect 219 18592 352 18598
rect 132 18550 138 18584
rect 172 18550 178 18584
rect 342 18582 352 18592
rect 858 18592 1619 18598
rect 858 18582 868 18592
rect 132 18392 178 18550
rect 970 18542 980 18552
rect 219 18536 980 18542
rect 1490 18542 1500 18552
rect 1490 18536 1619 18542
rect 219 18502 231 18536
rect 1607 18502 1619 18536
rect 219 18496 980 18502
rect 970 18486 980 18496
rect 1490 18496 1619 18502
rect 1490 18486 1500 18496
rect 1660 18488 1708 18646
rect 342 18446 352 18456
rect 219 18440 352 18446
rect 858 18446 868 18456
rect 1660 18454 1666 18488
rect 1700 18454 1708 18488
rect 858 18440 1619 18446
rect 219 18406 231 18440
rect 1607 18406 1619 18440
rect 219 18400 352 18406
rect 132 18358 138 18392
rect 172 18358 178 18392
rect 342 18390 352 18400
rect 858 18400 1619 18406
rect 858 18390 868 18400
rect 132 18200 178 18358
rect 970 18350 980 18360
rect 219 18344 980 18350
rect 1490 18350 1500 18360
rect 1490 18344 1619 18350
rect 219 18310 231 18344
rect 1607 18310 1619 18344
rect 219 18304 980 18310
rect 970 18294 980 18304
rect 1490 18304 1619 18310
rect 1490 18294 1500 18304
rect 1660 18296 1708 18454
rect 342 18254 352 18264
rect 219 18248 352 18254
rect 858 18254 868 18264
rect 1660 18262 1666 18296
rect 1700 18262 1708 18296
rect 858 18248 1619 18254
rect 219 18214 231 18248
rect 1607 18214 1619 18248
rect 219 18208 352 18214
rect 132 18166 138 18200
rect 172 18166 178 18200
rect 342 18198 352 18208
rect 858 18208 1619 18214
rect 858 18198 868 18208
rect 132 18008 178 18166
rect 970 18158 980 18168
rect 219 18152 980 18158
rect 1490 18158 1500 18168
rect 1490 18152 1619 18158
rect 219 18118 231 18152
rect 1607 18118 1619 18152
rect 219 18112 980 18118
rect 970 18102 980 18112
rect 1490 18112 1619 18118
rect 1490 18102 1500 18112
rect 1660 18104 1708 18262
rect 342 18062 352 18072
rect 219 18056 352 18062
rect 858 18062 868 18072
rect 1660 18070 1666 18104
rect 1700 18070 1708 18104
rect 858 18056 1619 18062
rect 219 18022 231 18056
rect 1607 18022 1619 18056
rect 219 18016 352 18022
rect 132 17974 138 18008
rect 172 17974 178 18008
rect 342 18006 352 18016
rect 858 18016 1619 18022
rect 858 18006 868 18016
rect 132 17816 178 17974
rect 970 17966 980 17976
rect 219 17960 980 17966
rect 1490 17966 1500 17976
rect 1490 17960 1619 17966
rect 219 17926 231 17960
rect 1607 17926 1619 17960
rect 219 17920 980 17926
rect 970 17910 980 17920
rect 1490 17920 1619 17926
rect 1490 17910 1500 17920
rect 1660 17912 1708 18070
rect 342 17870 352 17880
rect 219 17864 352 17870
rect 858 17870 868 17880
rect 1660 17878 1666 17912
rect 1700 17878 1708 17912
rect 858 17864 1619 17870
rect 219 17830 231 17864
rect 1607 17830 1619 17864
rect 219 17824 352 17830
rect 132 17782 138 17816
rect 172 17782 178 17816
rect 342 17814 352 17824
rect 858 17824 1619 17830
rect 858 17814 868 17824
rect 132 17624 178 17782
rect 970 17774 980 17784
rect 219 17768 980 17774
rect 1490 17774 1500 17784
rect 1490 17768 1619 17774
rect 219 17734 231 17768
rect 1607 17734 1619 17768
rect 219 17728 980 17734
rect 970 17718 980 17728
rect 1490 17728 1619 17734
rect 1490 17718 1500 17728
rect 1660 17720 1708 17878
rect 342 17678 352 17688
rect 219 17672 352 17678
rect 858 17678 868 17688
rect 1660 17686 1666 17720
rect 1700 17686 1708 17720
rect 858 17672 1619 17678
rect 219 17638 231 17672
rect 1607 17638 1619 17672
rect 219 17632 352 17638
rect 132 17590 138 17624
rect 172 17590 178 17624
rect 342 17622 352 17632
rect 858 17632 1619 17638
rect 858 17622 868 17632
rect 132 17432 178 17590
rect 970 17582 980 17592
rect 219 17576 980 17582
rect 1490 17582 1500 17592
rect 1490 17576 1619 17582
rect 219 17542 231 17576
rect 1607 17542 1619 17576
rect 219 17536 980 17542
rect 970 17526 980 17536
rect 1490 17536 1619 17542
rect 1490 17526 1500 17536
rect 1660 17528 1708 17686
rect 342 17486 352 17496
rect 219 17480 352 17486
rect 858 17486 868 17496
rect 1660 17494 1666 17528
rect 1700 17494 1708 17528
rect 858 17480 1619 17486
rect 219 17446 231 17480
rect 1607 17446 1619 17480
rect 219 17440 352 17446
rect 132 17398 138 17432
rect 172 17398 178 17432
rect 342 17430 352 17440
rect 858 17440 1619 17446
rect 858 17430 868 17440
rect 132 17240 178 17398
rect 970 17390 980 17400
rect 219 17384 980 17390
rect 1490 17390 1500 17400
rect 1490 17384 1619 17390
rect 219 17350 231 17384
rect 1607 17350 1619 17384
rect 219 17344 980 17350
rect 970 17334 980 17344
rect 1490 17344 1619 17350
rect 1490 17334 1500 17344
rect 1660 17336 1708 17494
rect 342 17294 352 17304
rect 219 17288 352 17294
rect 858 17294 868 17304
rect 1660 17302 1666 17336
rect 1700 17302 1708 17336
rect 858 17288 1619 17294
rect 219 17254 231 17288
rect 1607 17254 1619 17288
rect 219 17248 352 17254
rect 132 17206 138 17240
rect 172 17206 178 17240
rect 342 17238 352 17248
rect 858 17248 1619 17254
rect 858 17238 868 17248
rect 132 17048 178 17206
rect 970 17198 980 17208
rect 219 17192 980 17198
rect 1490 17198 1500 17208
rect 1490 17192 1619 17198
rect 219 17158 231 17192
rect 1607 17158 1619 17192
rect 219 17152 980 17158
rect 970 17142 980 17152
rect 1490 17152 1619 17158
rect 1490 17142 1500 17152
rect 1660 17144 1708 17302
rect 342 17102 352 17112
rect 219 17096 352 17102
rect 858 17102 868 17112
rect 1660 17110 1666 17144
rect 1700 17110 1708 17144
rect 858 17096 1619 17102
rect 219 17062 231 17096
rect 1607 17062 1619 17096
rect 219 17056 352 17062
rect 132 17014 138 17048
rect 172 17014 178 17048
rect 342 17046 352 17056
rect 858 17056 1619 17062
rect 858 17046 868 17056
rect 132 16856 178 17014
rect 970 17006 980 17016
rect 219 17000 980 17006
rect 1490 17006 1500 17016
rect 1490 17000 1619 17006
rect 219 16966 231 17000
rect 1607 16966 1619 17000
rect 219 16960 980 16966
rect 970 16950 980 16960
rect 1490 16960 1619 16966
rect 1490 16950 1500 16960
rect 1660 16952 1708 17110
rect 342 16910 352 16920
rect 219 16904 352 16910
rect 858 16910 868 16920
rect 1660 16918 1666 16952
rect 1700 16918 1708 16952
rect 858 16904 1619 16910
rect 219 16870 231 16904
rect 1607 16870 1619 16904
rect 219 16864 352 16870
rect 132 16822 138 16856
rect 172 16822 178 16856
rect 342 16854 352 16864
rect 858 16864 1619 16870
rect 858 16854 868 16864
rect 132 16664 178 16822
rect 970 16814 980 16824
rect 219 16808 980 16814
rect 1490 16814 1500 16824
rect 1490 16808 1619 16814
rect 219 16774 231 16808
rect 1607 16774 1619 16808
rect 219 16768 980 16774
rect 970 16758 980 16768
rect 1490 16768 1619 16774
rect 1490 16758 1500 16768
rect 1660 16760 1708 16918
rect 342 16718 352 16728
rect 219 16712 352 16718
rect 858 16718 868 16728
rect 1660 16726 1666 16760
rect 1700 16726 1708 16760
rect 858 16712 1619 16718
rect 219 16678 231 16712
rect 1607 16678 1619 16712
rect 219 16672 352 16678
rect 132 16630 138 16664
rect 172 16630 178 16664
rect 342 16662 352 16672
rect 858 16672 1619 16678
rect 858 16662 868 16672
rect 132 16472 178 16630
rect 970 16622 980 16632
rect 219 16616 980 16622
rect 1490 16622 1500 16632
rect 1490 16616 1619 16622
rect 219 16582 231 16616
rect 1607 16582 1619 16616
rect 219 16576 980 16582
rect 970 16566 980 16576
rect 1490 16576 1619 16582
rect 1490 16566 1500 16576
rect 1660 16568 1708 16726
rect 342 16526 352 16536
rect 219 16520 352 16526
rect 858 16526 868 16536
rect 1660 16534 1666 16568
rect 1700 16534 1708 16568
rect 858 16520 1619 16526
rect 219 16486 231 16520
rect 1607 16486 1619 16520
rect 219 16480 352 16486
rect 132 16438 138 16472
rect 172 16438 178 16472
rect 342 16470 352 16480
rect 858 16480 1619 16486
rect 858 16470 868 16480
rect 132 16280 178 16438
rect 970 16430 980 16440
rect 219 16424 980 16430
rect 1490 16430 1500 16440
rect 1490 16424 1619 16430
rect 219 16390 231 16424
rect 1607 16390 1619 16424
rect 219 16384 980 16390
rect 970 16374 980 16384
rect 1490 16384 1619 16390
rect 1490 16374 1500 16384
rect 1660 16376 1708 16534
rect 342 16334 352 16344
rect 219 16328 352 16334
rect 858 16334 868 16344
rect 1660 16342 1666 16376
rect 1700 16342 1708 16376
rect 858 16328 1619 16334
rect 219 16294 231 16328
rect 1607 16294 1619 16328
rect 219 16288 352 16294
rect 132 16246 138 16280
rect 172 16246 178 16280
rect 342 16278 352 16288
rect 858 16288 1619 16294
rect 858 16278 868 16288
rect 132 16088 178 16246
rect 970 16238 980 16248
rect 219 16232 980 16238
rect 1490 16238 1500 16248
rect 1490 16232 1619 16238
rect 219 16198 231 16232
rect 1607 16198 1619 16232
rect 219 16192 980 16198
rect 970 16182 980 16192
rect 1490 16192 1619 16198
rect 1490 16182 1500 16192
rect 1660 16184 1708 16342
rect 342 16142 352 16152
rect 219 16136 352 16142
rect 858 16142 868 16152
rect 1660 16150 1666 16184
rect 1700 16150 1708 16184
rect 858 16136 1619 16142
rect 219 16102 231 16136
rect 1607 16102 1619 16136
rect 219 16096 352 16102
rect 132 16054 138 16088
rect 172 16054 178 16088
rect 342 16086 352 16096
rect 858 16096 1619 16102
rect 858 16086 868 16096
rect 132 15896 178 16054
rect 970 16046 980 16056
rect 219 16040 980 16046
rect 1490 16046 1500 16056
rect 1490 16040 1619 16046
rect 219 16006 231 16040
rect 1607 16006 1619 16040
rect 219 16000 980 16006
rect 970 15990 980 16000
rect 1490 16000 1619 16006
rect 1490 15990 1500 16000
rect 1660 15992 1708 16150
rect 342 15950 352 15960
rect 219 15944 352 15950
rect 858 15950 868 15960
rect 1660 15958 1666 15992
rect 1700 15958 1708 15992
rect 858 15944 1619 15950
rect 219 15910 231 15944
rect 1607 15910 1619 15944
rect 219 15904 352 15910
rect 132 15862 138 15896
rect 172 15862 178 15896
rect 342 15894 352 15904
rect 858 15904 1619 15910
rect 858 15894 868 15904
rect 132 15704 178 15862
rect 970 15854 980 15864
rect 219 15848 980 15854
rect 1490 15854 1500 15864
rect 1490 15848 1619 15854
rect 219 15814 231 15848
rect 1607 15814 1619 15848
rect 219 15808 980 15814
rect 970 15798 980 15808
rect 1490 15808 1619 15814
rect 1490 15798 1500 15808
rect 1660 15800 1708 15958
rect 342 15758 352 15768
rect 219 15752 352 15758
rect 858 15758 868 15768
rect 1660 15766 1666 15800
rect 1700 15766 1708 15800
rect 858 15752 1619 15758
rect 219 15718 231 15752
rect 1607 15718 1619 15752
rect 219 15712 352 15718
rect 132 15670 138 15704
rect 172 15670 178 15704
rect 342 15702 352 15712
rect 858 15712 1619 15718
rect 858 15702 868 15712
rect 132 15512 178 15670
rect 970 15662 980 15672
rect 219 15656 980 15662
rect 1490 15662 1500 15672
rect 1490 15656 1619 15662
rect 219 15622 231 15656
rect 1607 15622 1619 15656
rect 219 15616 980 15622
rect 970 15606 980 15616
rect 1490 15616 1619 15622
rect 1490 15606 1500 15616
rect 1660 15608 1708 15766
rect 342 15566 352 15576
rect 219 15560 352 15566
rect 858 15566 868 15576
rect 1660 15574 1666 15608
rect 1700 15574 1708 15608
rect 858 15560 1619 15566
rect 219 15526 231 15560
rect 1607 15526 1619 15560
rect 219 15520 352 15526
rect 132 15478 138 15512
rect 172 15478 178 15512
rect 342 15510 352 15520
rect 858 15520 1619 15526
rect 858 15510 868 15520
rect 132 15320 178 15478
rect 970 15470 980 15480
rect 219 15464 980 15470
rect 1490 15470 1500 15480
rect 1490 15464 1619 15470
rect 219 15430 231 15464
rect 1607 15430 1619 15464
rect 219 15424 980 15430
rect 970 15414 980 15424
rect 1490 15424 1619 15430
rect 1490 15414 1500 15424
rect 1660 15416 1708 15574
rect 342 15374 352 15384
rect 219 15368 352 15374
rect 858 15374 868 15384
rect 1660 15382 1666 15416
rect 1700 15382 1708 15416
rect 858 15368 1619 15374
rect 219 15334 231 15368
rect 1607 15334 1619 15368
rect 219 15328 352 15334
rect 132 15286 138 15320
rect 172 15286 178 15320
rect 342 15318 352 15328
rect 858 15328 1619 15334
rect 858 15318 868 15328
rect 132 15128 178 15286
rect 970 15278 980 15288
rect 219 15272 980 15278
rect 1490 15278 1500 15288
rect 1490 15272 1619 15278
rect 219 15238 231 15272
rect 1607 15238 1619 15272
rect 219 15232 980 15238
rect 970 15222 980 15232
rect 1490 15232 1619 15238
rect 1490 15222 1500 15232
rect 1660 15224 1708 15382
rect 342 15182 352 15192
rect 219 15176 352 15182
rect 858 15182 868 15192
rect 1660 15190 1666 15224
rect 1700 15190 1708 15224
rect 858 15176 1619 15182
rect 219 15142 231 15176
rect 1607 15142 1619 15176
rect 219 15136 352 15142
rect 132 15094 138 15128
rect 172 15094 178 15128
rect 342 15126 352 15136
rect 858 15136 1619 15142
rect 858 15126 868 15136
rect 132 14936 178 15094
rect 970 15086 980 15096
rect 219 15080 980 15086
rect 1490 15086 1500 15096
rect 1490 15080 1619 15086
rect 219 15046 231 15080
rect 1607 15046 1619 15080
rect 219 15040 980 15046
rect 970 15030 980 15040
rect 1490 15040 1619 15046
rect 1490 15030 1500 15040
rect 1660 15032 1708 15190
rect 342 14990 352 15000
rect 219 14984 352 14990
rect 858 14990 868 15000
rect 1660 14998 1666 15032
rect 1700 14998 1708 15032
rect 858 14984 1619 14990
rect 219 14950 231 14984
rect 1607 14950 1619 14984
rect 219 14944 352 14950
rect 132 14902 138 14936
rect 172 14902 178 14936
rect 342 14934 352 14944
rect 858 14944 1619 14950
rect 858 14934 868 14944
rect 132 14744 178 14902
rect 970 14894 980 14904
rect 219 14888 980 14894
rect 1490 14894 1500 14904
rect 1490 14888 1619 14894
rect 219 14854 231 14888
rect 1607 14854 1619 14888
rect 219 14848 980 14854
rect 970 14838 980 14848
rect 1490 14848 1619 14854
rect 1490 14838 1500 14848
rect 1660 14840 1708 14998
rect 342 14798 352 14808
rect 219 14792 352 14798
rect 858 14798 868 14808
rect 1660 14806 1666 14840
rect 1700 14806 1708 14840
rect 858 14792 1619 14798
rect 219 14758 231 14792
rect 1607 14758 1619 14792
rect 219 14752 352 14758
rect 132 14710 138 14744
rect 172 14710 178 14744
rect 342 14742 352 14752
rect 858 14752 1619 14758
rect 858 14742 868 14752
rect 132 14552 178 14710
rect 970 14702 980 14712
rect 219 14696 980 14702
rect 1490 14702 1500 14712
rect 1490 14696 1619 14702
rect 219 14662 231 14696
rect 1607 14662 1619 14696
rect 219 14656 980 14662
rect 970 14646 980 14656
rect 1490 14656 1619 14662
rect 1490 14646 1500 14656
rect 1660 14648 1708 14806
rect 342 14606 352 14616
rect 219 14600 352 14606
rect 858 14606 868 14616
rect 1660 14614 1666 14648
rect 1700 14614 1708 14648
rect 858 14600 1619 14606
rect 219 14566 231 14600
rect 1607 14566 1619 14600
rect 219 14560 352 14566
rect 132 14518 138 14552
rect 172 14518 178 14552
rect 342 14550 352 14560
rect 858 14560 1619 14566
rect 858 14550 868 14560
rect 132 14360 178 14518
rect 970 14510 980 14520
rect 219 14504 980 14510
rect 1490 14510 1500 14520
rect 1490 14504 1619 14510
rect 219 14470 231 14504
rect 1607 14470 1619 14504
rect 219 14464 980 14470
rect 970 14454 980 14464
rect 1490 14464 1619 14470
rect 1490 14454 1500 14464
rect 1660 14456 1708 14614
rect 342 14414 352 14424
rect 219 14408 352 14414
rect 858 14414 868 14424
rect 1660 14422 1666 14456
rect 1700 14422 1708 14456
rect 858 14408 1619 14414
rect 219 14374 231 14408
rect 1607 14374 1619 14408
rect 219 14368 352 14374
rect 132 14326 138 14360
rect 172 14326 178 14360
rect 342 14358 352 14368
rect 858 14368 1619 14374
rect 858 14358 868 14368
rect 132 14168 178 14326
rect 970 14318 980 14328
rect 219 14312 980 14318
rect 1490 14318 1500 14328
rect 1490 14312 1619 14318
rect 219 14278 231 14312
rect 1607 14278 1619 14312
rect 219 14272 980 14278
rect 970 14262 980 14272
rect 1490 14272 1619 14278
rect 1490 14262 1500 14272
rect 1660 14264 1708 14422
rect 342 14222 352 14232
rect 219 14216 352 14222
rect 858 14222 868 14232
rect 1660 14230 1666 14264
rect 1700 14230 1708 14264
rect 858 14216 1619 14222
rect 219 14182 231 14216
rect 1607 14182 1619 14216
rect 219 14176 352 14182
rect 132 14134 138 14168
rect 172 14134 178 14168
rect 342 14166 352 14176
rect 858 14176 1619 14182
rect 858 14166 868 14176
rect 132 13976 178 14134
rect 970 14126 980 14136
rect 219 14120 980 14126
rect 1490 14126 1500 14136
rect 1490 14120 1619 14126
rect 219 14086 231 14120
rect 1607 14086 1619 14120
rect 219 14080 980 14086
rect 970 14070 980 14080
rect 1490 14080 1619 14086
rect 1490 14070 1500 14080
rect 1660 14072 1708 14230
rect 342 14030 352 14040
rect 219 14024 352 14030
rect 858 14030 868 14040
rect 1660 14038 1666 14072
rect 1700 14038 1708 14072
rect 858 14024 1619 14030
rect 219 13990 231 14024
rect 1607 13990 1619 14024
rect 219 13984 352 13990
rect 132 13942 138 13976
rect 172 13942 178 13976
rect 342 13974 352 13984
rect 858 13984 1619 13990
rect 858 13974 868 13984
rect 132 13784 178 13942
rect 970 13934 980 13944
rect 219 13928 980 13934
rect 1490 13934 1500 13944
rect 1490 13928 1619 13934
rect 219 13894 231 13928
rect 1607 13894 1619 13928
rect 219 13888 980 13894
rect 970 13878 980 13888
rect 1490 13888 1619 13894
rect 1490 13878 1500 13888
rect 1660 13880 1708 14038
rect 342 13838 352 13848
rect 219 13832 352 13838
rect 858 13838 868 13848
rect 1660 13846 1666 13880
rect 1700 13846 1708 13880
rect 858 13832 1619 13838
rect 219 13798 231 13832
rect 1607 13798 1619 13832
rect 219 13792 352 13798
rect 132 13750 138 13784
rect 172 13750 178 13784
rect 342 13782 352 13792
rect 858 13792 1619 13798
rect 858 13782 868 13792
rect 132 13592 178 13750
rect 970 13742 980 13752
rect 219 13736 980 13742
rect 1490 13742 1500 13752
rect 1490 13736 1619 13742
rect 219 13702 231 13736
rect 1607 13702 1619 13736
rect 219 13696 980 13702
rect 970 13686 980 13696
rect 1490 13696 1619 13702
rect 1490 13686 1500 13696
rect 1660 13688 1708 13846
rect 342 13646 352 13656
rect 219 13640 352 13646
rect 858 13646 868 13656
rect 1660 13654 1666 13688
rect 1700 13654 1708 13688
rect 858 13640 1619 13646
rect 219 13606 231 13640
rect 1607 13606 1619 13640
rect 219 13600 352 13606
rect 132 13558 138 13592
rect 172 13558 178 13592
rect 342 13590 352 13600
rect 858 13600 1619 13606
rect 858 13590 868 13600
rect 132 13400 178 13558
rect 970 13550 980 13560
rect 219 13544 980 13550
rect 1490 13550 1500 13560
rect 1490 13544 1619 13550
rect 219 13510 231 13544
rect 1607 13510 1619 13544
rect 219 13504 980 13510
rect 970 13494 980 13504
rect 1490 13504 1619 13510
rect 1490 13494 1500 13504
rect 1660 13496 1708 13654
rect 342 13454 352 13464
rect 219 13448 352 13454
rect 858 13454 868 13464
rect 1660 13462 1666 13496
rect 1700 13462 1708 13496
rect 858 13448 1619 13454
rect 219 13414 231 13448
rect 1607 13414 1619 13448
rect 219 13408 352 13414
rect 132 13366 138 13400
rect 172 13366 178 13400
rect 342 13398 352 13408
rect 858 13408 1619 13414
rect 858 13398 868 13408
rect 132 13208 178 13366
rect 970 13358 980 13368
rect 219 13352 980 13358
rect 1490 13358 1500 13368
rect 1490 13352 1619 13358
rect 219 13318 231 13352
rect 1607 13318 1619 13352
rect 219 13312 980 13318
rect 970 13302 980 13312
rect 1490 13312 1619 13318
rect 1490 13302 1500 13312
rect 1660 13304 1708 13462
rect 342 13262 352 13272
rect 219 13256 352 13262
rect 858 13262 868 13272
rect 1660 13270 1666 13304
rect 1700 13270 1708 13304
rect 858 13256 1619 13262
rect 219 13222 231 13256
rect 1607 13222 1619 13256
rect 219 13216 352 13222
rect 132 13174 138 13208
rect 172 13174 178 13208
rect 342 13206 352 13216
rect 858 13216 1619 13222
rect 858 13206 868 13216
rect 132 13016 178 13174
rect 970 13166 980 13176
rect 219 13160 980 13166
rect 1490 13166 1500 13176
rect 1490 13160 1619 13166
rect 219 13126 231 13160
rect 1607 13126 1619 13160
rect 219 13120 980 13126
rect 970 13110 980 13120
rect 1490 13120 1619 13126
rect 1490 13110 1500 13120
rect 1660 13112 1708 13270
rect 342 13070 352 13080
rect 219 13064 352 13070
rect 858 13070 868 13080
rect 1660 13078 1666 13112
rect 1700 13078 1708 13112
rect 858 13064 1619 13070
rect 219 13030 231 13064
rect 1607 13030 1619 13064
rect 219 13024 352 13030
rect 132 12982 138 13016
rect 172 12982 178 13016
rect 342 13014 352 13024
rect 858 13024 1619 13030
rect 858 13014 868 13024
rect 132 12824 178 12982
rect 970 12974 980 12984
rect 219 12968 980 12974
rect 1490 12974 1500 12984
rect 1490 12968 1619 12974
rect 219 12934 231 12968
rect 1607 12934 1619 12968
rect 219 12928 980 12934
rect 970 12918 980 12928
rect 1490 12928 1619 12934
rect 1490 12918 1500 12928
rect 1660 12920 1708 13078
rect 342 12878 352 12888
rect 219 12872 352 12878
rect 858 12878 868 12888
rect 1660 12886 1666 12920
rect 1700 12886 1708 12920
rect 858 12872 1619 12878
rect 219 12838 231 12872
rect 1607 12838 1619 12872
rect 219 12832 352 12838
rect 132 12790 138 12824
rect 172 12790 178 12824
rect 342 12822 352 12832
rect 858 12832 1619 12838
rect 858 12822 868 12832
rect 132 12632 178 12790
rect 970 12782 980 12792
rect 219 12776 980 12782
rect 1490 12782 1500 12792
rect 1490 12776 1619 12782
rect 219 12742 231 12776
rect 1607 12742 1619 12776
rect 219 12736 980 12742
rect 970 12726 980 12736
rect 1490 12736 1619 12742
rect 1490 12726 1500 12736
rect 1660 12728 1708 12886
rect 342 12686 352 12696
rect 219 12680 352 12686
rect 858 12686 868 12696
rect 1660 12694 1666 12728
rect 1700 12694 1708 12728
rect 858 12680 1619 12686
rect 219 12646 231 12680
rect 1607 12646 1619 12680
rect 219 12640 352 12646
rect 132 12598 138 12632
rect 172 12598 178 12632
rect 342 12630 352 12640
rect 858 12640 1619 12646
rect 858 12630 868 12640
rect 132 12440 178 12598
rect 970 12590 980 12600
rect 219 12584 980 12590
rect 1490 12590 1500 12600
rect 1490 12584 1619 12590
rect 219 12550 231 12584
rect 1607 12550 1619 12584
rect 219 12544 980 12550
rect 970 12534 980 12544
rect 1490 12544 1619 12550
rect 1490 12534 1500 12544
rect 1660 12536 1708 12694
rect 342 12494 352 12504
rect 219 12488 352 12494
rect 858 12494 868 12504
rect 1660 12502 1666 12536
rect 1700 12502 1708 12536
rect 858 12488 1619 12494
rect 219 12454 231 12488
rect 1607 12454 1619 12488
rect 219 12448 352 12454
rect 132 12406 138 12440
rect 172 12406 178 12440
rect 342 12438 352 12448
rect 858 12448 1619 12454
rect 858 12438 868 12448
rect 132 12248 178 12406
rect 970 12398 980 12408
rect 219 12392 980 12398
rect 1490 12398 1500 12408
rect 1490 12392 1619 12398
rect 219 12358 231 12392
rect 1607 12358 1619 12392
rect 219 12352 980 12358
rect 970 12342 980 12352
rect 1490 12352 1619 12358
rect 1490 12342 1500 12352
rect 1660 12344 1708 12502
rect 342 12302 352 12312
rect 219 12296 352 12302
rect 858 12302 868 12312
rect 1660 12310 1666 12344
rect 1700 12310 1708 12344
rect 858 12296 1619 12302
rect 219 12262 231 12296
rect 1607 12262 1619 12296
rect 219 12256 352 12262
rect 132 12214 138 12248
rect 172 12214 178 12248
rect 342 12246 352 12256
rect 858 12256 1619 12262
rect 858 12246 868 12256
rect 132 12056 178 12214
rect 970 12206 980 12216
rect 219 12200 980 12206
rect 1490 12206 1500 12216
rect 1490 12200 1619 12206
rect 219 12166 231 12200
rect 1607 12166 1619 12200
rect 219 12160 980 12166
rect 970 12150 980 12160
rect 1490 12160 1619 12166
rect 1490 12150 1500 12160
rect 1660 12152 1708 12310
rect 342 12110 352 12120
rect 219 12104 352 12110
rect 858 12110 868 12120
rect 1660 12118 1666 12152
rect 1700 12118 1708 12152
rect 858 12104 1619 12110
rect 219 12070 231 12104
rect 1607 12070 1619 12104
rect 219 12064 352 12070
rect 132 12022 138 12056
rect 172 12022 178 12056
rect 342 12054 352 12064
rect 858 12064 1619 12070
rect 858 12054 868 12064
rect 132 11864 178 12022
rect 970 12014 980 12024
rect 219 12008 980 12014
rect 1490 12014 1500 12024
rect 1490 12008 1619 12014
rect 219 11974 231 12008
rect 1607 11974 1619 12008
rect 219 11968 980 11974
rect 970 11958 980 11968
rect 1490 11968 1619 11974
rect 1490 11958 1500 11968
rect 1660 11960 1708 12118
rect 342 11918 352 11928
rect 219 11912 352 11918
rect 858 11918 868 11928
rect 1660 11926 1666 11960
rect 1700 11926 1708 11960
rect 858 11912 1619 11918
rect 219 11878 231 11912
rect 1607 11878 1619 11912
rect 219 11872 352 11878
rect 132 11830 138 11864
rect 172 11830 178 11864
rect 342 11862 352 11872
rect 858 11872 1619 11878
rect 858 11862 868 11872
rect 132 11672 178 11830
rect 970 11822 980 11832
rect 219 11816 980 11822
rect 1490 11822 1500 11832
rect 1490 11816 1619 11822
rect 219 11782 231 11816
rect 1607 11782 1619 11816
rect 219 11776 980 11782
rect 970 11766 980 11776
rect 1490 11776 1619 11782
rect 1490 11766 1500 11776
rect 1660 11768 1708 11926
rect 342 11726 352 11736
rect 219 11720 352 11726
rect 858 11726 868 11736
rect 1660 11734 1666 11768
rect 1700 11734 1708 11768
rect 858 11720 1619 11726
rect 219 11686 231 11720
rect 1607 11686 1619 11720
rect 219 11680 352 11686
rect 132 11638 138 11672
rect 172 11638 178 11672
rect 342 11670 352 11680
rect 858 11680 1619 11686
rect 858 11670 868 11680
rect 132 11480 178 11638
rect 970 11630 980 11640
rect 219 11624 980 11630
rect 1490 11630 1500 11640
rect 1490 11624 1619 11630
rect 219 11590 231 11624
rect 1607 11590 1619 11624
rect 219 11584 980 11590
rect 970 11574 980 11584
rect 1490 11584 1619 11590
rect 1490 11574 1500 11584
rect 1660 11576 1708 11734
rect 342 11534 352 11544
rect 219 11528 352 11534
rect 858 11534 868 11544
rect 1660 11542 1666 11576
rect 1700 11542 1708 11576
rect 858 11528 1619 11534
rect 219 11494 231 11528
rect 1607 11494 1619 11528
rect 219 11488 352 11494
rect 132 11446 138 11480
rect 172 11446 178 11480
rect 342 11478 352 11488
rect 858 11488 1619 11494
rect 858 11478 868 11488
rect 132 11288 178 11446
rect 970 11438 980 11448
rect 219 11432 980 11438
rect 1490 11438 1500 11448
rect 1490 11432 1619 11438
rect 219 11398 231 11432
rect 1607 11398 1619 11432
rect 219 11392 980 11398
rect 970 11382 980 11392
rect 1490 11392 1619 11398
rect 1490 11382 1500 11392
rect 1660 11384 1708 11542
rect 342 11342 352 11352
rect 219 11336 352 11342
rect 858 11342 868 11352
rect 1660 11350 1666 11384
rect 1700 11350 1708 11384
rect 858 11336 1619 11342
rect 219 11302 231 11336
rect 1607 11302 1619 11336
rect 219 11296 352 11302
rect 132 11254 138 11288
rect 172 11254 178 11288
rect 342 11286 352 11296
rect 858 11296 1619 11302
rect 858 11286 868 11296
rect 132 11096 178 11254
rect 970 11246 980 11256
rect 219 11240 980 11246
rect 1490 11246 1500 11256
rect 1490 11240 1619 11246
rect 219 11206 231 11240
rect 1607 11206 1619 11240
rect 219 11200 980 11206
rect 970 11190 980 11200
rect 1490 11200 1619 11206
rect 1490 11190 1500 11200
rect 1660 11192 1708 11350
rect 342 11150 352 11160
rect 219 11144 352 11150
rect 858 11150 868 11160
rect 1660 11158 1666 11192
rect 1700 11158 1708 11192
rect 858 11144 1619 11150
rect 219 11110 231 11144
rect 1607 11110 1619 11144
rect 219 11104 352 11110
rect 132 11062 138 11096
rect 172 11062 178 11096
rect 342 11094 352 11104
rect 858 11104 1619 11110
rect 858 11094 868 11104
rect 132 10904 178 11062
rect 970 11054 980 11064
rect 219 11048 980 11054
rect 1490 11054 1500 11064
rect 1490 11048 1619 11054
rect 219 11014 231 11048
rect 1607 11014 1619 11048
rect 219 11008 980 11014
rect 970 10998 980 11008
rect 1490 11008 1619 11014
rect 1490 10998 1500 11008
rect 1660 11000 1708 11158
rect 342 10958 352 10968
rect 219 10952 352 10958
rect 858 10958 868 10968
rect 1660 10966 1666 11000
rect 1700 10966 1708 11000
rect 858 10952 1619 10958
rect 219 10918 231 10952
rect 1607 10918 1619 10952
rect 219 10912 352 10918
rect 132 10870 138 10904
rect 172 10870 178 10904
rect 342 10902 352 10912
rect 858 10912 1619 10918
rect 858 10902 868 10912
rect 132 10712 178 10870
rect 970 10862 980 10872
rect 219 10856 980 10862
rect 1490 10862 1500 10872
rect 1490 10856 1619 10862
rect 219 10822 231 10856
rect 1607 10822 1619 10856
rect 219 10816 980 10822
rect 970 10806 980 10816
rect 1490 10816 1619 10822
rect 1490 10806 1500 10816
rect 1660 10808 1708 10966
rect 342 10766 352 10776
rect 219 10760 352 10766
rect 858 10766 868 10776
rect 1660 10774 1666 10808
rect 1700 10774 1708 10808
rect 858 10760 1619 10766
rect 219 10726 231 10760
rect 1607 10726 1619 10760
rect 219 10720 352 10726
rect 132 10678 138 10712
rect 172 10678 178 10712
rect 342 10710 352 10720
rect 858 10720 1619 10726
rect 858 10710 868 10720
rect 132 10520 178 10678
rect 970 10670 980 10680
rect 219 10664 980 10670
rect 1490 10670 1500 10680
rect 1490 10664 1619 10670
rect 219 10630 231 10664
rect 1607 10630 1619 10664
rect 219 10624 980 10630
rect 970 10614 980 10624
rect 1490 10624 1619 10630
rect 1490 10614 1500 10624
rect 1660 10616 1708 10774
rect 342 10574 352 10584
rect 219 10568 352 10574
rect 858 10574 868 10584
rect 1660 10582 1666 10616
rect 1700 10582 1708 10616
rect 858 10568 1619 10574
rect 219 10534 231 10568
rect 1607 10534 1619 10568
rect 219 10528 352 10534
rect 132 10486 138 10520
rect 172 10486 178 10520
rect 342 10518 352 10528
rect 858 10528 1619 10534
rect 858 10518 868 10528
rect 132 10328 178 10486
rect 970 10478 980 10488
rect 219 10472 980 10478
rect 1490 10478 1500 10488
rect 1490 10472 1619 10478
rect 219 10438 231 10472
rect 1607 10438 1619 10472
rect 219 10432 980 10438
rect 970 10422 980 10432
rect 1490 10432 1619 10438
rect 1490 10422 1500 10432
rect 1660 10424 1708 10582
rect 342 10382 352 10392
rect 219 10376 352 10382
rect 858 10382 868 10392
rect 1660 10390 1666 10424
rect 1700 10390 1708 10424
rect 858 10376 1619 10382
rect 219 10342 231 10376
rect 1607 10342 1619 10376
rect 219 10336 352 10342
rect 132 10294 138 10328
rect 172 10294 178 10328
rect 342 10326 352 10336
rect 858 10336 1619 10342
rect 858 10326 868 10336
rect 132 10136 178 10294
rect 970 10286 980 10296
rect 219 10280 980 10286
rect 1490 10286 1500 10296
rect 1490 10280 1619 10286
rect 219 10246 231 10280
rect 1607 10246 1619 10280
rect 219 10240 980 10246
rect 970 10230 980 10240
rect 1490 10240 1619 10246
rect 1490 10230 1500 10240
rect 1660 10232 1708 10390
rect 342 10190 352 10200
rect 219 10184 352 10190
rect 858 10190 868 10200
rect 1660 10198 1666 10232
rect 1700 10198 1708 10232
rect 858 10184 1619 10190
rect 219 10150 231 10184
rect 1607 10150 1619 10184
rect 219 10144 352 10150
rect 132 10102 138 10136
rect 172 10102 178 10136
rect 342 10134 352 10144
rect 858 10144 1619 10150
rect 858 10134 868 10144
rect 132 9944 178 10102
rect 970 10094 980 10104
rect 219 10088 980 10094
rect 1490 10094 1500 10104
rect 1490 10088 1619 10094
rect 219 10054 231 10088
rect 1607 10054 1619 10088
rect 219 10048 980 10054
rect 970 10038 980 10048
rect 1490 10048 1619 10054
rect 1490 10038 1500 10048
rect 1660 10040 1708 10198
rect 342 9998 352 10008
rect 219 9992 352 9998
rect 858 9998 868 10008
rect 1660 10006 1666 10040
rect 1700 10006 1708 10040
rect 858 9992 1619 9998
rect 219 9958 231 9992
rect 1607 9958 1619 9992
rect 219 9952 352 9958
rect 132 9910 138 9944
rect 172 9910 178 9944
rect 342 9942 352 9952
rect 858 9952 1619 9958
rect 858 9942 868 9952
rect 132 9752 178 9910
rect 970 9902 980 9912
rect 219 9896 980 9902
rect 1490 9902 1500 9912
rect 1490 9896 1619 9902
rect 219 9862 231 9896
rect 1607 9862 1619 9896
rect 219 9856 980 9862
rect 970 9846 980 9856
rect 1490 9856 1619 9862
rect 1490 9846 1500 9856
rect 1660 9848 1708 10006
rect 342 9806 352 9816
rect 219 9800 352 9806
rect 858 9806 868 9816
rect 1660 9814 1666 9848
rect 1700 9814 1708 9848
rect 858 9800 1619 9806
rect 219 9766 231 9800
rect 1607 9766 1619 9800
rect 219 9760 352 9766
rect 132 9718 138 9752
rect 172 9718 178 9752
rect 342 9750 352 9760
rect 858 9760 1619 9766
rect 858 9750 868 9760
rect 132 9560 178 9718
rect 970 9710 980 9720
rect 219 9704 980 9710
rect 1490 9710 1500 9720
rect 1490 9704 1619 9710
rect 219 9670 231 9704
rect 1607 9670 1619 9704
rect 219 9664 980 9670
rect 970 9654 980 9664
rect 1490 9664 1619 9670
rect 1490 9654 1500 9664
rect 1660 9656 1708 9814
rect 342 9614 352 9624
rect 219 9608 352 9614
rect 858 9614 868 9624
rect 1660 9622 1666 9656
rect 1700 9622 1708 9656
rect 858 9608 1619 9614
rect 219 9574 231 9608
rect 1607 9574 1619 9608
rect 219 9568 352 9574
rect 132 9526 138 9560
rect 172 9526 178 9560
rect 342 9558 352 9568
rect 858 9568 1619 9574
rect 858 9558 868 9568
rect 132 9368 178 9526
rect 970 9518 980 9528
rect 219 9512 980 9518
rect 1490 9518 1500 9528
rect 1490 9512 1619 9518
rect 219 9478 231 9512
rect 1607 9478 1619 9512
rect 219 9472 980 9478
rect 970 9462 980 9472
rect 1490 9472 1619 9478
rect 1490 9462 1500 9472
rect 1660 9464 1708 9622
rect 342 9422 352 9432
rect 219 9416 352 9422
rect 858 9422 868 9432
rect 1660 9430 1666 9464
rect 1700 9430 1708 9464
rect 858 9416 1619 9422
rect 219 9382 231 9416
rect 1607 9382 1619 9416
rect 219 9376 352 9382
rect 132 9334 138 9368
rect 172 9334 178 9368
rect 342 9366 352 9376
rect 858 9376 1619 9382
rect 858 9366 868 9376
rect 132 9176 178 9334
rect 970 9326 980 9336
rect 219 9320 980 9326
rect 1490 9326 1500 9336
rect 1490 9320 1619 9326
rect 219 9286 231 9320
rect 1607 9286 1619 9320
rect 219 9280 980 9286
rect 970 9270 980 9280
rect 1490 9280 1619 9286
rect 1490 9270 1500 9280
rect 1660 9272 1708 9430
rect 342 9230 352 9240
rect 219 9224 352 9230
rect 858 9230 868 9240
rect 1660 9238 1666 9272
rect 1700 9238 1708 9272
rect 858 9224 1619 9230
rect 219 9190 231 9224
rect 1607 9190 1619 9224
rect 219 9184 352 9190
rect 132 9142 138 9176
rect 172 9142 178 9176
rect 342 9174 352 9184
rect 858 9184 1619 9190
rect 858 9174 868 9184
rect 132 8984 178 9142
rect 970 9134 980 9144
rect 219 9128 980 9134
rect 1490 9134 1500 9144
rect 1490 9128 1619 9134
rect 219 9094 231 9128
rect 1607 9094 1619 9128
rect 219 9088 980 9094
rect 970 9078 980 9088
rect 1490 9088 1619 9094
rect 1490 9078 1500 9088
rect 1660 9080 1708 9238
rect 342 9038 352 9048
rect 219 9032 352 9038
rect 858 9038 868 9048
rect 1660 9046 1666 9080
rect 1700 9046 1708 9080
rect 858 9032 1619 9038
rect 219 8998 231 9032
rect 1607 8998 1619 9032
rect 219 8992 352 8998
rect 132 8950 138 8984
rect 172 8950 178 8984
rect 342 8982 352 8992
rect 858 8992 1619 8998
rect 858 8982 868 8992
rect 132 8792 178 8950
rect 970 8942 980 8952
rect 219 8936 980 8942
rect 1490 8942 1500 8952
rect 1490 8936 1619 8942
rect 219 8902 231 8936
rect 1607 8902 1619 8936
rect 219 8896 980 8902
rect 970 8886 980 8896
rect 1490 8896 1619 8902
rect 1490 8886 1500 8896
rect 1660 8888 1708 9046
rect 342 8846 352 8856
rect 219 8840 352 8846
rect 858 8846 868 8856
rect 1660 8854 1666 8888
rect 1700 8854 1708 8888
rect 858 8840 1619 8846
rect 219 8806 231 8840
rect 1607 8806 1619 8840
rect 219 8800 352 8806
rect 132 8758 138 8792
rect 172 8758 178 8792
rect 342 8790 352 8800
rect 858 8800 1619 8806
rect 858 8790 868 8800
rect 132 8600 178 8758
rect 970 8750 980 8760
rect 219 8744 980 8750
rect 1490 8750 1500 8760
rect 1490 8744 1619 8750
rect 219 8710 231 8744
rect 1607 8710 1619 8744
rect 219 8704 980 8710
rect 970 8694 980 8704
rect 1490 8704 1619 8710
rect 1490 8694 1500 8704
rect 1660 8696 1708 8854
rect 342 8654 352 8664
rect 219 8648 352 8654
rect 858 8654 868 8664
rect 1660 8662 1666 8696
rect 1700 8662 1708 8696
rect 858 8648 1619 8654
rect 219 8614 231 8648
rect 1607 8614 1619 8648
rect 219 8608 352 8614
rect 132 8566 138 8600
rect 172 8566 178 8600
rect 342 8598 352 8608
rect 858 8608 1619 8614
rect 858 8598 868 8608
rect 132 8408 178 8566
rect 970 8558 980 8568
rect 219 8552 980 8558
rect 1490 8558 1500 8568
rect 1490 8552 1619 8558
rect 219 8518 231 8552
rect 1607 8518 1619 8552
rect 219 8512 980 8518
rect 970 8502 980 8512
rect 1490 8512 1619 8518
rect 1490 8502 1500 8512
rect 1660 8504 1708 8662
rect 342 8462 352 8472
rect 219 8456 352 8462
rect 858 8462 868 8472
rect 1660 8470 1666 8504
rect 1700 8470 1708 8504
rect 858 8456 1619 8462
rect 219 8422 231 8456
rect 1607 8422 1619 8456
rect 219 8416 352 8422
rect 132 8374 138 8408
rect 172 8374 178 8408
rect 342 8406 352 8416
rect 858 8416 1619 8422
rect 858 8406 868 8416
rect 132 8216 178 8374
rect 970 8366 980 8376
rect 219 8360 980 8366
rect 1490 8366 1500 8376
rect 1490 8360 1619 8366
rect 219 8326 231 8360
rect 1607 8326 1619 8360
rect 219 8320 980 8326
rect 970 8310 980 8320
rect 1490 8320 1619 8326
rect 1490 8310 1500 8320
rect 1660 8312 1708 8470
rect 342 8270 352 8280
rect 219 8264 352 8270
rect 858 8270 868 8280
rect 1660 8278 1666 8312
rect 1700 8278 1708 8312
rect 858 8264 1619 8270
rect 219 8230 231 8264
rect 1607 8230 1619 8264
rect 219 8224 352 8230
rect 132 8182 138 8216
rect 172 8182 178 8216
rect 342 8214 352 8224
rect 858 8224 1619 8230
rect 858 8214 868 8224
rect 132 8024 178 8182
rect 970 8174 980 8184
rect 219 8168 980 8174
rect 1490 8174 1500 8184
rect 1490 8168 1619 8174
rect 219 8134 231 8168
rect 1607 8134 1619 8168
rect 219 8128 980 8134
rect 970 8118 980 8128
rect 1490 8128 1619 8134
rect 1490 8118 1500 8128
rect 1660 8120 1708 8278
rect 342 8078 352 8088
rect 219 8072 352 8078
rect 858 8078 868 8088
rect 1660 8086 1666 8120
rect 1700 8086 1708 8120
rect 858 8072 1619 8078
rect 219 8038 231 8072
rect 1607 8038 1619 8072
rect 219 8032 352 8038
rect 132 7990 138 8024
rect 172 7990 178 8024
rect 342 8022 352 8032
rect 858 8032 1619 8038
rect 858 8022 868 8032
rect 132 7832 178 7990
rect 970 7982 980 7992
rect 219 7976 980 7982
rect 1490 7982 1500 7992
rect 1490 7976 1619 7982
rect 219 7942 231 7976
rect 1607 7942 1619 7976
rect 219 7936 980 7942
rect 970 7926 980 7936
rect 1490 7936 1619 7942
rect 1490 7926 1500 7936
rect 1660 7928 1708 8086
rect 342 7886 352 7896
rect 219 7880 352 7886
rect 858 7886 868 7896
rect 1660 7894 1666 7928
rect 1700 7894 1708 7928
rect 858 7880 1619 7886
rect 219 7846 231 7880
rect 1607 7846 1619 7880
rect 219 7840 352 7846
rect 132 7798 138 7832
rect 172 7798 178 7832
rect 342 7830 352 7840
rect 858 7840 1619 7846
rect 858 7830 868 7840
rect 132 7640 178 7798
rect 970 7790 980 7800
rect 219 7784 980 7790
rect 1490 7790 1500 7800
rect 1490 7784 1619 7790
rect 219 7750 231 7784
rect 1607 7750 1619 7784
rect 219 7744 980 7750
rect 970 7734 980 7744
rect 1490 7744 1619 7750
rect 1490 7734 1500 7744
rect 1660 7736 1708 7894
rect 342 7694 352 7704
rect 219 7688 352 7694
rect 858 7694 868 7704
rect 1660 7702 1666 7736
rect 1700 7702 1708 7736
rect 858 7688 1619 7694
rect 219 7654 231 7688
rect 1607 7654 1619 7688
rect 219 7648 352 7654
rect 132 7606 138 7640
rect 172 7606 178 7640
rect 342 7638 352 7648
rect 858 7648 1619 7654
rect 858 7638 868 7648
rect 132 7448 178 7606
rect 970 7598 980 7608
rect 219 7592 980 7598
rect 1490 7598 1500 7608
rect 1490 7592 1619 7598
rect 219 7558 231 7592
rect 1607 7558 1619 7592
rect 219 7552 980 7558
rect 970 7542 980 7552
rect 1490 7552 1619 7558
rect 1490 7542 1500 7552
rect 1660 7544 1708 7702
rect 342 7502 352 7512
rect 219 7496 352 7502
rect 858 7502 868 7512
rect 1660 7510 1666 7544
rect 1700 7510 1708 7544
rect 858 7496 1619 7502
rect 219 7462 231 7496
rect 1607 7462 1619 7496
rect 219 7456 352 7462
rect 132 7414 138 7448
rect 172 7414 178 7448
rect 342 7446 352 7456
rect 858 7456 1619 7462
rect 858 7446 868 7456
rect 132 7256 178 7414
rect 970 7406 980 7416
rect 219 7400 980 7406
rect 1490 7406 1500 7416
rect 1490 7400 1619 7406
rect 219 7366 231 7400
rect 1607 7366 1619 7400
rect 219 7360 980 7366
rect 970 7350 980 7360
rect 1490 7360 1619 7366
rect 1490 7350 1500 7360
rect 1660 7352 1708 7510
rect 342 7310 352 7320
rect 219 7304 352 7310
rect 858 7310 868 7320
rect 1660 7318 1666 7352
rect 1700 7318 1708 7352
rect 858 7304 1619 7310
rect 219 7270 231 7304
rect 1607 7270 1619 7304
rect 219 7264 352 7270
rect 132 7222 138 7256
rect 172 7222 178 7256
rect 342 7254 352 7264
rect 858 7264 1619 7270
rect 858 7254 868 7264
rect 132 7064 178 7222
rect 970 7214 980 7224
rect 219 7208 980 7214
rect 1490 7214 1500 7224
rect 1490 7208 1619 7214
rect 219 7174 231 7208
rect 1607 7174 1619 7208
rect 219 7168 980 7174
rect 970 7158 980 7168
rect 1490 7168 1619 7174
rect 1490 7158 1500 7168
rect 1660 7160 1708 7318
rect 342 7118 352 7128
rect 219 7112 352 7118
rect 858 7118 868 7128
rect 1660 7126 1666 7160
rect 1700 7126 1708 7160
rect 858 7112 1619 7118
rect 219 7078 231 7112
rect 1607 7078 1619 7112
rect 219 7072 352 7078
rect 132 7030 138 7064
rect 172 7030 178 7064
rect 342 7062 352 7072
rect 858 7072 1619 7078
rect 858 7062 868 7072
rect 132 6872 178 7030
rect 970 7022 980 7032
rect 219 7016 980 7022
rect 1490 7022 1500 7032
rect 1490 7016 1619 7022
rect 219 6982 231 7016
rect 1607 6982 1619 7016
rect 219 6976 980 6982
rect 970 6966 980 6976
rect 1490 6976 1619 6982
rect 1490 6966 1500 6976
rect 1660 6968 1708 7126
rect 342 6926 352 6936
rect 219 6920 352 6926
rect 858 6926 868 6936
rect 1660 6934 1666 6968
rect 1700 6934 1708 6968
rect 858 6920 1619 6926
rect 219 6886 231 6920
rect 1607 6886 1619 6920
rect 219 6880 352 6886
rect 132 6838 138 6872
rect 172 6838 178 6872
rect 342 6870 352 6880
rect 858 6880 1619 6886
rect 858 6870 868 6880
rect 132 6680 178 6838
rect 970 6830 980 6840
rect 219 6824 980 6830
rect 1490 6830 1500 6840
rect 1490 6824 1619 6830
rect 219 6790 231 6824
rect 1607 6790 1619 6824
rect 219 6784 980 6790
rect 970 6774 980 6784
rect 1490 6784 1619 6790
rect 1490 6774 1500 6784
rect 1660 6776 1708 6934
rect 342 6734 352 6744
rect 219 6728 352 6734
rect 858 6734 868 6744
rect 1660 6742 1666 6776
rect 1700 6742 1708 6776
rect 858 6728 1619 6734
rect 219 6694 231 6728
rect 1607 6694 1619 6728
rect 219 6688 352 6694
rect 132 6646 138 6680
rect 172 6646 178 6680
rect 342 6678 352 6688
rect 858 6688 1619 6694
rect 858 6678 868 6688
rect 132 6488 178 6646
rect 970 6638 980 6648
rect 219 6632 980 6638
rect 1490 6638 1500 6648
rect 1490 6632 1619 6638
rect 219 6598 231 6632
rect 1607 6598 1619 6632
rect 219 6592 980 6598
rect 970 6582 980 6592
rect 1490 6592 1619 6598
rect 1490 6582 1500 6592
rect 1660 6584 1708 6742
rect 342 6542 352 6552
rect 219 6536 352 6542
rect 858 6542 868 6552
rect 1660 6550 1666 6584
rect 1700 6550 1708 6584
rect 858 6536 1619 6542
rect 219 6502 231 6536
rect 1607 6502 1619 6536
rect 219 6496 352 6502
rect 132 6454 138 6488
rect 172 6454 178 6488
rect 342 6486 352 6496
rect 858 6496 1619 6502
rect 858 6486 868 6496
rect 132 6296 178 6454
rect 970 6446 980 6456
rect 219 6440 980 6446
rect 1490 6446 1500 6456
rect 1490 6440 1619 6446
rect 219 6406 231 6440
rect 1607 6406 1619 6440
rect 219 6400 980 6406
rect 970 6390 980 6400
rect 1490 6400 1619 6406
rect 1490 6390 1500 6400
rect 1660 6392 1708 6550
rect 342 6350 352 6360
rect 219 6344 352 6350
rect 858 6350 868 6360
rect 1660 6358 1666 6392
rect 1700 6358 1708 6392
rect 858 6344 1619 6350
rect 219 6310 231 6344
rect 1607 6310 1619 6344
rect 219 6304 352 6310
rect 132 6262 138 6296
rect 172 6262 178 6296
rect 342 6294 352 6304
rect 858 6304 1619 6310
rect 858 6294 868 6304
rect 132 6104 178 6262
rect 970 6254 980 6264
rect 219 6248 980 6254
rect 1490 6254 1500 6264
rect 1490 6248 1619 6254
rect 219 6214 231 6248
rect 1607 6214 1619 6248
rect 219 6208 980 6214
rect 970 6198 980 6208
rect 1490 6208 1619 6214
rect 1490 6198 1500 6208
rect 1660 6200 1708 6358
rect 342 6158 352 6168
rect 219 6152 352 6158
rect 858 6158 868 6168
rect 1660 6166 1666 6200
rect 1700 6166 1708 6200
rect 858 6152 1619 6158
rect 219 6118 231 6152
rect 1607 6118 1619 6152
rect 219 6112 352 6118
rect 132 6070 138 6104
rect 172 6070 178 6104
rect 342 6102 352 6112
rect 858 6112 1619 6118
rect 858 6102 868 6112
rect 132 5912 178 6070
rect 970 6062 980 6072
rect 219 6056 980 6062
rect 1490 6062 1500 6072
rect 1490 6056 1619 6062
rect 219 6022 231 6056
rect 1607 6022 1619 6056
rect 219 6016 980 6022
rect 970 6006 980 6016
rect 1490 6016 1619 6022
rect 1490 6006 1500 6016
rect 1660 6008 1708 6166
rect 342 5966 352 5976
rect 219 5960 352 5966
rect 858 5966 868 5976
rect 1660 5974 1666 6008
rect 1700 5974 1708 6008
rect 858 5960 1619 5966
rect 219 5926 231 5960
rect 1607 5926 1619 5960
rect 219 5920 352 5926
rect 132 5878 138 5912
rect 172 5878 178 5912
rect 342 5910 352 5920
rect 858 5920 1619 5926
rect 858 5910 868 5920
rect 132 5720 178 5878
rect 970 5870 980 5880
rect 219 5864 980 5870
rect 1490 5870 1500 5880
rect 1490 5864 1619 5870
rect 219 5830 231 5864
rect 1607 5830 1619 5864
rect 219 5824 980 5830
rect 970 5814 980 5824
rect 1490 5824 1619 5830
rect 1490 5814 1500 5824
rect 1660 5816 1708 5974
rect 342 5774 352 5784
rect 219 5768 352 5774
rect 858 5774 868 5784
rect 1660 5782 1666 5816
rect 1700 5782 1708 5816
rect 858 5768 1619 5774
rect 219 5734 231 5768
rect 1607 5734 1619 5768
rect 219 5728 352 5734
rect 132 5686 138 5720
rect 172 5686 178 5720
rect 342 5718 352 5728
rect 858 5728 1619 5734
rect 858 5718 868 5728
rect 132 5528 178 5686
rect 970 5678 980 5688
rect 219 5672 980 5678
rect 1490 5678 1500 5688
rect 1490 5672 1619 5678
rect 219 5638 231 5672
rect 1607 5638 1619 5672
rect 219 5632 980 5638
rect 970 5622 980 5632
rect 1490 5632 1619 5638
rect 1490 5622 1500 5632
rect 1660 5624 1708 5782
rect 342 5582 352 5592
rect 219 5576 352 5582
rect 858 5582 868 5592
rect 1660 5590 1666 5624
rect 1700 5590 1708 5624
rect 858 5576 1619 5582
rect 219 5542 231 5576
rect 1607 5542 1619 5576
rect 219 5536 352 5542
rect 132 5494 138 5528
rect 172 5494 178 5528
rect 342 5526 352 5536
rect 858 5536 1619 5542
rect 858 5526 868 5536
rect 132 5336 178 5494
rect 970 5486 980 5496
rect 219 5480 980 5486
rect 1490 5486 1500 5496
rect 1490 5480 1619 5486
rect 219 5446 231 5480
rect 1607 5446 1619 5480
rect 219 5440 980 5446
rect 970 5430 980 5440
rect 1490 5440 1619 5446
rect 1490 5430 1500 5440
rect 1660 5432 1708 5590
rect 342 5390 352 5400
rect 219 5384 352 5390
rect 858 5390 868 5400
rect 1660 5398 1666 5432
rect 1700 5398 1708 5432
rect 858 5384 1619 5390
rect 219 5350 231 5384
rect 1607 5350 1619 5384
rect 219 5344 352 5350
rect 132 5302 138 5336
rect 172 5302 178 5336
rect 342 5334 352 5344
rect 858 5344 1619 5350
rect 858 5334 868 5344
rect 132 5144 178 5302
rect 970 5294 980 5304
rect 219 5288 980 5294
rect 1490 5294 1500 5304
rect 1490 5288 1619 5294
rect 219 5254 231 5288
rect 1607 5254 1619 5288
rect 219 5248 980 5254
rect 970 5238 980 5248
rect 1490 5248 1619 5254
rect 1490 5238 1500 5248
rect 1660 5240 1708 5398
rect 342 5198 352 5208
rect 219 5192 352 5198
rect 858 5198 868 5208
rect 1660 5206 1666 5240
rect 1700 5206 1708 5240
rect 858 5192 1619 5198
rect 219 5158 231 5192
rect 1607 5158 1619 5192
rect 219 5152 352 5158
rect 132 5110 138 5144
rect 172 5110 178 5144
rect 342 5142 352 5152
rect 858 5152 1619 5158
rect 858 5142 868 5152
rect 132 4952 178 5110
rect 970 5102 980 5112
rect 219 5096 980 5102
rect 1490 5102 1500 5112
rect 1490 5096 1619 5102
rect 219 5062 231 5096
rect 1607 5062 1619 5096
rect 219 5056 980 5062
rect 970 5046 980 5056
rect 1490 5056 1619 5062
rect 1490 5046 1500 5056
rect 1660 5048 1708 5206
rect 342 5006 352 5016
rect 219 5000 352 5006
rect 858 5006 868 5016
rect 1660 5014 1666 5048
rect 1700 5014 1708 5048
rect 858 5000 1619 5006
rect 219 4966 231 5000
rect 1607 4966 1619 5000
rect 219 4960 352 4966
rect 132 4918 138 4952
rect 172 4918 178 4952
rect 342 4950 352 4960
rect 858 4960 1619 4966
rect 858 4950 868 4960
rect 132 4760 178 4918
rect 970 4910 980 4920
rect 219 4904 980 4910
rect 1490 4910 1500 4920
rect 1490 4904 1619 4910
rect 219 4870 231 4904
rect 1607 4870 1619 4904
rect 219 4864 980 4870
rect 970 4854 980 4864
rect 1490 4864 1619 4870
rect 1490 4854 1500 4864
rect 1660 4856 1708 5014
rect 342 4814 352 4824
rect 219 4808 352 4814
rect 858 4814 868 4824
rect 1660 4822 1666 4856
rect 1700 4822 1708 4856
rect 858 4808 1619 4814
rect 219 4774 231 4808
rect 1607 4774 1619 4808
rect 219 4768 352 4774
rect 132 4726 138 4760
rect 172 4726 178 4760
rect 342 4758 352 4768
rect 858 4768 1619 4774
rect 858 4758 868 4768
rect 132 4568 178 4726
rect 970 4718 980 4728
rect 219 4712 980 4718
rect 1490 4718 1500 4728
rect 1490 4712 1619 4718
rect 219 4678 231 4712
rect 1607 4678 1619 4712
rect 219 4672 980 4678
rect 970 4662 980 4672
rect 1490 4672 1619 4678
rect 1490 4662 1500 4672
rect 1660 4664 1708 4822
rect 342 4622 352 4632
rect 219 4616 352 4622
rect 858 4622 868 4632
rect 1660 4630 1666 4664
rect 1700 4630 1708 4664
rect 858 4616 1619 4622
rect 219 4582 231 4616
rect 1607 4582 1619 4616
rect 219 4576 352 4582
rect 132 4534 138 4568
rect 172 4534 178 4568
rect 342 4566 352 4576
rect 858 4576 1619 4582
rect 858 4566 868 4576
rect 132 4376 178 4534
rect 970 4526 980 4536
rect 219 4520 980 4526
rect 1490 4526 1500 4536
rect 1490 4520 1619 4526
rect 219 4486 231 4520
rect 1607 4486 1619 4520
rect 219 4480 980 4486
rect 970 4470 980 4480
rect 1490 4480 1619 4486
rect 1490 4470 1500 4480
rect 1660 4472 1708 4630
rect 342 4430 352 4440
rect 219 4424 352 4430
rect 858 4430 868 4440
rect 1660 4438 1666 4472
rect 1700 4438 1708 4472
rect 858 4424 1619 4430
rect 219 4390 231 4424
rect 1607 4390 1619 4424
rect 219 4384 352 4390
rect 132 4342 138 4376
rect 172 4342 178 4376
rect 342 4374 352 4384
rect 858 4384 1619 4390
rect 858 4374 868 4384
rect 132 4184 178 4342
rect 970 4334 980 4344
rect 219 4328 980 4334
rect 1490 4334 1500 4344
rect 1490 4328 1619 4334
rect 219 4294 231 4328
rect 1607 4294 1619 4328
rect 219 4288 980 4294
rect 970 4278 980 4288
rect 1490 4288 1619 4294
rect 1490 4278 1500 4288
rect 1660 4280 1708 4438
rect 342 4238 352 4248
rect 219 4232 352 4238
rect 858 4238 868 4248
rect 1660 4246 1666 4280
rect 1700 4246 1708 4280
rect 858 4232 1619 4238
rect 219 4198 231 4232
rect 1607 4198 1619 4232
rect 219 4192 352 4198
rect 132 4150 138 4184
rect 172 4150 178 4184
rect 342 4182 352 4192
rect 858 4192 1619 4198
rect 858 4182 868 4192
rect 132 3992 178 4150
rect 970 4142 980 4152
rect 219 4136 980 4142
rect 1490 4142 1500 4152
rect 1490 4136 1619 4142
rect 219 4102 231 4136
rect 1607 4102 1619 4136
rect 219 4096 980 4102
rect 970 4086 980 4096
rect 1490 4096 1619 4102
rect 1490 4086 1500 4096
rect 1660 4088 1708 4246
rect 342 4046 352 4056
rect 219 4040 352 4046
rect 858 4046 868 4056
rect 1660 4054 1666 4088
rect 1700 4054 1708 4088
rect 858 4040 1619 4046
rect 219 4006 231 4040
rect 1607 4006 1619 4040
rect 219 4000 352 4006
rect 132 3958 138 3992
rect 172 3958 178 3992
rect 342 3990 352 4000
rect 858 4000 1619 4006
rect 858 3990 868 4000
rect 132 3800 178 3958
rect 970 3950 980 3960
rect 219 3944 980 3950
rect 1490 3950 1500 3960
rect 1490 3944 1619 3950
rect 219 3910 231 3944
rect 1607 3910 1619 3944
rect 219 3904 980 3910
rect 970 3894 980 3904
rect 1490 3904 1619 3910
rect 1490 3894 1500 3904
rect 1660 3896 1708 4054
rect 342 3854 352 3864
rect 219 3848 352 3854
rect 858 3854 868 3864
rect 1660 3862 1666 3896
rect 1700 3862 1708 3896
rect 858 3848 1619 3854
rect 219 3814 231 3848
rect 1607 3814 1619 3848
rect 219 3808 352 3814
rect 132 3766 138 3800
rect 172 3766 178 3800
rect 342 3798 352 3808
rect 858 3808 1619 3814
rect 858 3798 868 3808
rect 132 3608 178 3766
rect 970 3758 980 3768
rect 219 3752 980 3758
rect 1490 3758 1500 3768
rect 1490 3752 1619 3758
rect 219 3718 231 3752
rect 1607 3718 1619 3752
rect 219 3712 980 3718
rect 970 3702 980 3712
rect 1490 3712 1619 3718
rect 1490 3702 1500 3712
rect 1660 3704 1708 3862
rect 342 3662 352 3672
rect 219 3656 352 3662
rect 858 3662 868 3672
rect 1660 3670 1666 3704
rect 1700 3670 1708 3704
rect 858 3656 1619 3662
rect 219 3622 231 3656
rect 1607 3622 1619 3656
rect 219 3616 352 3622
rect 132 3574 138 3608
rect 172 3574 178 3608
rect 342 3606 352 3616
rect 858 3616 1619 3622
rect 858 3606 868 3616
rect 132 3416 178 3574
rect 970 3566 980 3576
rect 219 3560 980 3566
rect 1490 3566 1500 3576
rect 1490 3560 1619 3566
rect 219 3526 231 3560
rect 1607 3526 1619 3560
rect 219 3520 980 3526
rect 970 3510 980 3520
rect 1490 3520 1619 3526
rect 1490 3510 1500 3520
rect 1660 3512 1708 3670
rect 342 3470 352 3480
rect 219 3464 352 3470
rect 858 3470 868 3480
rect 1660 3478 1666 3512
rect 1700 3478 1708 3512
rect 858 3464 1619 3470
rect 219 3430 231 3464
rect 1607 3430 1619 3464
rect 219 3424 352 3430
rect 132 3382 138 3416
rect 172 3382 178 3416
rect 342 3414 352 3424
rect 858 3424 1619 3430
rect 858 3414 868 3424
rect 132 3224 178 3382
rect 970 3374 980 3384
rect 219 3368 980 3374
rect 1490 3374 1500 3384
rect 1490 3368 1619 3374
rect 219 3334 231 3368
rect 1607 3334 1619 3368
rect 219 3328 980 3334
rect 970 3318 980 3328
rect 1490 3328 1619 3334
rect 1490 3318 1500 3328
rect 1660 3320 1708 3478
rect 342 3278 352 3288
rect 219 3272 352 3278
rect 858 3278 868 3288
rect 1660 3286 1666 3320
rect 1700 3286 1708 3320
rect 858 3272 1619 3278
rect 219 3238 231 3272
rect 1607 3238 1619 3272
rect 219 3232 352 3238
rect 132 3190 138 3224
rect 172 3190 178 3224
rect 342 3222 352 3232
rect 858 3232 1619 3238
rect 858 3222 868 3232
rect 132 3032 178 3190
rect 970 3182 980 3192
rect 219 3176 980 3182
rect 1490 3182 1500 3192
rect 1490 3176 1619 3182
rect 219 3142 231 3176
rect 1607 3142 1619 3176
rect 219 3136 980 3142
rect 970 3126 980 3136
rect 1490 3136 1619 3142
rect 1490 3126 1500 3136
rect 1660 3128 1708 3286
rect 342 3086 352 3096
rect 219 3080 352 3086
rect 858 3086 868 3096
rect 1660 3094 1666 3128
rect 1700 3094 1708 3128
rect 858 3080 1619 3086
rect 219 3046 231 3080
rect 1607 3046 1619 3080
rect 219 3040 352 3046
rect 132 2998 138 3032
rect 172 2998 178 3032
rect 342 3030 352 3040
rect 858 3040 1619 3046
rect 858 3030 868 3040
rect 132 2840 178 2998
rect 970 2990 980 3000
rect 219 2984 980 2990
rect 1490 2990 1500 3000
rect 1490 2984 1619 2990
rect 219 2950 231 2984
rect 1607 2950 1619 2984
rect 219 2944 980 2950
rect 970 2934 980 2944
rect 1490 2944 1619 2950
rect 1490 2934 1500 2944
rect 1660 2936 1708 3094
rect 342 2894 352 2904
rect 219 2888 352 2894
rect 858 2894 868 2904
rect 1660 2902 1666 2936
rect 1700 2902 1708 2936
rect 858 2888 1619 2894
rect 219 2854 231 2888
rect 1607 2854 1619 2888
rect 219 2848 352 2854
rect 132 2806 138 2840
rect 172 2806 178 2840
rect 342 2838 352 2848
rect 858 2848 1619 2854
rect 858 2838 868 2848
rect 132 2648 178 2806
rect 970 2798 980 2808
rect 219 2792 980 2798
rect 1490 2798 1500 2808
rect 1490 2792 1619 2798
rect 219 2758 231 2792
rect 1607 2758 1619 2792
rect 219 2752 980 2758
rect 970 2742 980 2752
rect 1490 2752 1619 2758
rect 1490 2742 1500 2752
rect 1660 2744 1708 2902
rect 342 2702 352 2712
rect 219 2696 352 2702
rect 858 2702 868 2712
rect 1660 2710 1666 2744
rect 1700 2710 1708 2744
rect 858 2696 1619 2702
rect 219 2662 231 2696
rect 1607 2662 1619 2696
rect 219 2656 352 2662
rect 132 2614 138 2648
rect 172 2614 178 2648
rect 342 2646 352 2656
rect 858 2656 1619 2662
rect 858 2646 868 2656
rect 132 2456 178 2614
rect 970 2606 980 2616
rect 219 2600 980 2606
rect 1490 2606 1500 2616
rect 1490 2600 1619 2606
rect 219 2566 231 2600
rect 1607 2566 1619 2600
rect 219 2560 980 2566
rect 970 2550 980 2560
rect 1490 2560 1619 2566
rect 1490 2550 1500 2560
rect 1660 2552 1708 2710
rect 342 2510 352 2520
rect 219 2504 352 2510
rect 858 2510 868 2520
rect 1660 2518 1666 2552
rect 1700 2518 1708 2552
rect 858 2504 1619 2510
rect 219 2470 231 2504
rect 1607 2470 1619 2504
rect 219 2464 352 2470
rect 132 2422 138 2456
rect 172 2422 178 2456
rect 342 2454 352 2464
rect 858 2464 1619 2470
rect 858 2454 868 2464
rect 132 2264 178 2422
rect 970 2414 980 2424
rect 219 2408 980 2414
rect 1490 2414 1500 2424
rect 1490 2408 1619 2414
rect 219 2374 231 2408
rect 1607 2374 1619 2408
rect 219 2368 980 2374
rect 970 2358 980 2368
rect 1490 2368 1619 2374
rect 1490 2358 1500 2368
rect 1660 2360 1708 2518
rect 342 2318 352 2328
rect 219 2312 352 2318
rect 858 2318 868 2328
rect 1660 2326 1666 2360
rect 1700 2326 1708 2360
rect 858 2312 1619 2318
rect 219 2278 231 2312
rect 1607 2278 1619 2312
rect 219 2272 352 2278
rect 132 2230 138 2264
rect 172 2230 178 2264
rect 342 2262 352 2272
rect 858 2272 1619 2278
rect 858 2262 868 2272
rect 132 2072 178 2230
rect 970 2222 980 2232
rect 219 2216 980 2222
rect 1490 2222 1500 2232
rect 1490 2216 1619 2222
rect 219 2182 231 2216
rect 1607 2182 1619 2216
rect 219 2176 980 2182
rect 970 2166 980 2176
rect 1490 2176 1619 2182
rect 1490 2166 1500 2176
rect 1660 2168 1708 2326
rect 342 2126 352 2136
rect 219 2120 352 2126
rect 858 2126 868 2136
rect 1660 2134 1666 2168
rect 1700 2134 1708 2168
rect 858 2120 1619 2126
rect 219 2086 231 2120
rect 1607 2086 1619 2120
rect 219 2080 352 2086
rect 132 2038 138 2072
rect 172 2038 178 2072
rect 342 2070 352 2080
rect 858 2080 1619 2086
rect 858 2070 868 2080
rect 132 1880 178 2038
rect 970 2030 980 2040
rect 219 2024 980 2030
rect 1490 2030 1500 2040
rect 1490 2024 1619 2030
rect 219 1990 231 2024
rect 1607 1990 1619 2024
rect 219 1984 980 1990
rect 970 1974 980 1984
rect 1490 1984 1619 1990
rect 1490 1974 1500 1984
rect 1660 1976 1708 2134
rect 342 1934 352 1944
rect 219 1928 352 1934
rect 858 1934 868 1944
rect 1660 1942 1666 1976
rect 1700 1942 1708 1976
rect 858 1928 1619 1934
rect 219 1894 231 1928
rect 1607 1894 1619 1928
rect 219 1888 352 1894
rect 132 1846 138 1880
rect 172 1846 178 1880
rect 342 1878 352 1888
rect 858 1888 1619 1894
rect 858 1878 868 1888
rect 132 1688 178 1846
rect 970 1838 980 1848
rect 219 1832 980 1838
rect 1490 1838 1500 1848
rect 1490 1832 1619 1838
rect 219 1798 231 1832
rect 1607 1798 1619 1832
rect 219 1792 980 1798
rect 970 1782 980 1792
rect 1490 1792 1619 1798
rect 1490 1782 1500 1792
rect 1660 1784 1708 1942
rect 342 1742 352 1752
rect 219 1736 352 1742
rect 858 1742 868 1752
rect 1660 1750 1666 1784
rect 1700 1750 1708 1784
rect 858 1736 1619 1742
rect 219 1702 231 1736
rect 1607 1702 1619 1736
rect 219 1696 352 1702
rect 132 1654 138 1688
rect 172 1654 178 1688
rect 342 1686 352 1696
rect 858 1696 1619 1702
rect 858 1686 868 1696
rect 132 1496 178 1654
rect 970 1646 980 1656
rect 219 1640 980 1646
rect 1490 1646 1500 1656
rect 1490 1640 1619 1646
rect 219 1606 231 1640
rect 1607 1606 1619 1640
rect 219 1600 980 1606
rect 970 1590 980 1600
rect 1490 1600 1619 1606
rect 1490 1590 1500 1600
rect 1660 1592 1708 1750
rect 342 1550 352 1560
rect 219 1544 352 1550
rect 858 1550 868 1560
rect 1660 1558 1666 1592
rect 1700 1558 1708 1592
rect 858 1544 1619 1550
rect 219 1510 231 1544
rect 1607 1510 1619 1544
rect 219 1504 352 1510
rect 132 1462 138 1496
rect 172 1462 178 1496
rect 342 1494 352 1504
rect 858 1504 1619 1510
rect 858 1494 868 1504
rect 132 1304 178 1462
rect 970 1454 980 1464
rect 219 1448 980 1454
rect 1490 1454 1500 1464
rect 1490 1448 1619 1454
rect 219 1414 231 1448
rect 1607 1414 1619 1448
rect 219 1408 980 1414
rect 970 1398 980 1408
rect 1490 1408 1619 1414
rect 1490 1398 1500 1408
rect 1660 1400 1708 1558
rect 342 1358 352 1368
rect 219 1352 352 1358
rect 858 1358 868 1368
rect 1660 1366 1666 1400
rect 1700 1366 1708 1400
rect 858 1352 1619 1358
rect 219 1318 231 1352
rect 1607 1318 1619 1352
rect 219 1312 352 1318
rect 132 1270 138 1304
rect 172 1270 178 1304
rect 342 1302 352 1312
rect 858 1312 1619 1318
rect 858 1302 868 1312
rect 132 1112 178 1270
rect 970 1262 980 1272
rect 219 1256 980 1262
rect 1490 1262 1500 1272
rect 1490 1256 1619 1262
rect 219 1222 231 1256
rect 1607 1222 1619 1256
rect 219 1216 980 1222
rect 970 1206 980 1216
rect 1490 1216 1619 1222
rect 1490 1206 1500 1216
rect 1660 1208 1708 1366
rect 342 1166 352 1176
rect 219 1160 352 1166
rect 858 1166 868 1176
rect 1660 1174 1666 1208
rect 1700 1174 1708 1208
rect 858 1160 1619 1166
rect 219 1126 231 1160
rect 1607 1126 1619 1160
rect 219 1120 352 1126
rect 132 1078 138 1112
rect 172 1078 178 1112
rect 342 1110 352 1120
rect 858 1120 1619 1126
rect 858 1110 868 1120
rect 132 920 178 1078
rect 970 1070 980 1080
rect 219 1064 980 1070
rect 1490 1070 1500 1080
rect 1490 1064 1619 1070
rect 219 1030 231 1064
rect 1607 1030 1619 1064
rect 219 1024 980 1030
rect 970 1014 980 1024
rect 1490 1024 1619 1030
rect 1490 1014 1500 1024
rect 1660 1016 1708 1174
rect 342 974 352 984
rect 219 968 352 974
rect 858 974 868 984
rect 1660 982 1666 1016
rect 1700 982 1708 1016
rect 858 968 1619 974
rect 219 934 231 968
rect 1607 934 1619 968
rect 219 928 352 934
rect 132 886 138 920
rect 172 886 178 920
rect 342 918 352 928
rect 858 928 1619 934
rect 858 918 868 928
rect 132 728 178 886
rect 970 878 980 888
rect 219 872 980 878
rect 1490 878 1500 888
rect 1490 872 1619 878
rect 219 838 231 872
rect 1607 838 1619 872
rect 219 832 980 838
rect 970 822 980 832
rect 1490 832 1619 838
rect 1490 822 1500 832
rect 1660 824 1708 982
rect 342 782 352 792
rect 219 776 352 782
rect 858 782 868 792
rect 1660 790 1666 824
rect 1700 790 1708 824
rect 858 776 1619 782
rect 219 742 231 776
rect 1607 742 1619 776
rect 219 736 352 742
rect 132 694 138 728
rect 172 694 178 728
rect 342 726 352 736
rect 858 736 1619 742
rect 858 726 868 736
rect 132 682 178 694
rect 970 686 980 696
rect 219 680 980 686
rect 1490 686 1500 696
rect 1490 680 1619 686
rect 219 646 231 680
rect 1607 646 1619 680
rect 219 640 980 646
rect 970 630 980 640
rect 1490 640 1619 646
rect 1490 630 1500 640
rect 1660 632 1708 790
rect 342 590 352 600
rect 219 584 352 590
rect 858 590 868 600
rect 1660 598 1666 632
rect 1700 598 1706 632
rect 858 584 1619 590
rect 1660 584 1706 598
rect 219 550 231 584
rect 1607 550 1619 584
rect 219 544 352 550
rect 342 534 352 544
rect 858 544 1619 550
rect 858 534 868 544
<< via1 >>
rect 132 45072 1706 45126
rect 352 44202 858 44218
rect 352 44168 858 44202
rect 352 44152 858 44168
rect 980 44106 1490 44122
rect 980 44072 1490 44106
rect 980 44056 1490 44072
rect 352 44010 858 44026
rect 352 43976 858 44010
rect 352 43960 858 43976
rect 980 43914 1490 43930
rect 980 43880 1490 43914
rect 980 43864 1490 43880
rect 352 43818 858 43834
rect 352 43784 858 43818
rect 352 43768 858 43784
rect 980 43722 1490 43738
rect 980 43688 1490 43722
rect 980 43672 1490 43688
rect 352 43626 858 43642
rect 352 43592 858 43626
rect 352 43576 858 43592
rect 980 43530 1490 43546
rect 980 43496 1490 43530
rect 980 43480 1490 43496
rect 352 43434 858 43450
rect 352 43400 858 43434
rect 352 43384 858 43400
rect 980 43338 1490 43354
rect 980 43304 1490 43338
rect 980 43288 1490 43304
rect 352 43242 858 43258
rect 352 43208 858 43242
rect 352 43192 858 43208
rect 980 43146 1490 43162
rect 980 43112 1490 43146
rect 980 43096 1490 43112
rect 352 43050 858 43066
rect 352 43016 858 43050
rect 352 43000 858 43016
rect 980 42954 1490 42970
rect 980 42920 1490 42954
rect 980 42904 1490 42920
rect 352 42858 858 42874
rect 352 42824 858 42858
rect 352 42808 858 42824
rect 980 42762 1490 42778
rect 980 42728 1490 42762
rect 980 42712 1490 42728
rect 352 42666 858 42682
rect 352 42632 858 42666
rect 352 42616 858 42632
rect 980 42570 1490 42586
rect 980 42536 1490 42570
rect 980 42520 1490 42536
rect 352 42474 858 42490
rect 352 42440 858 42474
rect 352 42424 858 42440
rect 980 42378 1490 42394
rect 980 42344 1490 42378
rect 980 42328 1490 42344
rect 352 42282 858 42298
rect 352 42248 858 42282
rect 352 42232 858 42248
rect 980 42186 1490 42202
rect 980 42152 1490 42186
rect 980 42136 1490 42152
rect 352 42090 858 42106
rect 352 42056 858 42090
rect 352 42040 858 42056
rect 980 41994 1490 42010
rect 980 41960 1490 41994
rect 980 41944 1490 41960
rect 352 41898 858 41914
rect 352 41864 858 41898
rect 352 41848 858 41864
rect 980 41802 1490 41818
rect 980 41768 1490 41802
rect 980 41752 1490 41768
rect 352 41706 858 41722
rect 352 41672 858 41706
rect 352 41656 858 41672
rect 980 41610 1490 41626
rect 980 41576 1490 41610
rect 980 41560 1490 41576
rect 352 41514 858 41530
rect 352 41480 858 41514
rect 352 41464 858 41480
rect 980 41418 1490 41434
rect 980 41384 1490 41418
rect 980 41368 1490 41384
rect 352 41322 858 41338
rect 352 41288 858 41322
rect 352 41272 858 41288
rect 980 41226 1490 41242
rect 980 41192 1490 41226
rect 980 41176 1490 41192
rect 352 41130 858 41146
rect 352 41096 858 41130
rect 352 41080 858 41096
rect 980 41034 1490 41050
rect 980 41000 1490 41034
rect 980 40984 1490 41000
rect 352 40938 858 40954
rect 352 40904 858 40938
rect 352 40888 858 40904
rect 980 40842 1490 40858
rect 980 40808 1490 40842
rect 980 40792 1490 40808
rect 352 40746 858 40762
rect 352 40712 858 40746
rect 352 40696 858 40712
rect 980 40650 1490 40666
rect 980 40616 1490 40650
rect 980 40600 1490 40616
rect 352 40554 858 40570
rect 352 40520 858 40554
rect 352 40504 858 40520
rect 980 40458 1490 40474
rect 980 40424 1490 40458
rect 980 40408 1490 40424
rect 352 40362 858 40378
rect 352 40328 858 40362
rect 352 40312 858 40328
rect 980 40266 1490 40282
rect 980 40232 1490 40266
rect 980 40216 1490 40232
rect 352 40170 858 40186
rect 352 40136 858 40170
rect 352 40120 858 40136
rect 980 40074 1490 40090
rect 980 40040 1490 40074
rect 980 40024 1490 40040
rect 352 39978 858 39994
rect 352 39944 858 39978
rect 352 39928 858 39944
rect 980 39882 1490 39898
rect 980 39848 1490 39882
rect 980 39832 1490 39848
rect 352 39786 858 39802
rect 352 39752 858 39786
rect 352 39736 858 39752
rect 980 39690 1490 39706
rect 980 39656 1490 39690
rect 980 39640 1490 39656
rect 352 39594 858 39610
rect 352 39560 858 39594
rect 352 39544 858 39560
rect 980 39498 1490 39514
rect 980 39464 1490 39498
rect 980 39448 1490 39464
rect 352 39402 858 39418
rect 352 39368 858 39402
rect 352 39352 858 39368
rect 980 39306 1490 39322
rect 980 39272 1490 39306
rect 980 39256 1490 39272
rect 352 39210 858 39226
rect 352 39176 858 39210
rect 352 39160 858 39176
rect 980 39114 1490 39130
rect 980 39080 1490 39114
rect 980 39064 1490 39080
rect 352 39018 858 39034
rect 352 38984 858 39018
rect 352 38968 858 38984
rect 980 38922 1490 38938
rect 980 38888 1490 38922
rect 980 38872 1490 38888
rect 352 38826 858 38842
rect 352 38792 858 38826
rect 352 38776 858 38792
rect 980 38730 1490 38746
rect 980 38696 1490 38730
rect 980 38680 1490 38696
rect 352 38634 858 38650
rect 352 38600 858 38634
rect 352 38584 858 38600
rect 980 38538 1490 38554
rect 980 38504 1490 38538
rect 980 38488 1490 38504
rect 352 38442 858 38458
rect 352 38408 858 38442
rect 352 38392 858 38408
rect 980 38346 1490 38362
rect 980 38312 1490 38346
rect 980 38296 1490 38312
rect 352 38250 858 38266
rect 352 38216 858 38250
rect 352 38200 858 38216
rect 980 38154 1490 38170
rect 980 38120 1490 38154
rect 980 38104 1490 38120
rect 352 38058 858 38074
rect 352 38024 858 38058
rect 352 38008 858 38024
rect 980 37962 1490 37978
rect 980 37928 1490 37962
rect 980 37912 1490 37928
rect 352 37866 858 37882
rect 352 37832 858 37866
rect 352 37816 858 37832
rect 980 37770 1490 37786
rect 980 37736 1490 37770
rect 980 37720 1490 37736
rect 352 37674 858 37690
rect 352 37640 858 37674
rect 352 37624 858 37640
rect 980 37578 1490 37594
rect 980 37544 1490 37578
rect 980 37528 1490 37544
rect 352 37482 858 37498
rect 352 37448 858 37482
rect 352 37432 858 37448
rect 980 37386 1490 37402
rect 980 37352 1490 37386
rect 980 37336 1490 37352
rect 352 37290 858 37306
rect 352 37256 858 37290
rect 352 37240 858 37256
rect 980 37194 1490 37210
rect 980 37160 1490 37194
rect 980 37144 1490 37160
rect 352 37098 858 37114
rect 352 37064 858 37098
rect 352 37048 858 37064
rect 980 37002 1490 37018
rect 980 36968 1490 37002
rect 980 36952 1490 36968
rect 352 36906 858 36922
rect 352 36872 858 36906
rect 352 36856 858 36872
rect 980 36810 1490 36826
rect 980 36776 1490 36810
rect 980 36760 1490 36776
rect 352 36714 858 36730
rect 352 36680 858 36714
rect 352 36664 858 36680
rect 980 36618 1490 36634
rect 980 36584 1490 36618
rect 980 36568 1490 36584
rect 352 36522 858 36538
rect 352 36488 858 36522
rect 352 36472 858 36488
rect 980 36426 1490 36442
rect 980 36392 1490 36426
rect 980 36376 1490 36392
rect 352 36330 858 36346
rect 352 36296 858 36330
rect 352 36280 858 36296
rect 980 36234 1490 36250
rect 980 36200 1490 36234
rect 980 36184 1490 36200
rect 352 36138 858 36154
rect 352 36104 858 36138
rect 352 36088 858 36104
rect 980 36042 1490 36058
rect 980 36008 1490 36042
rect 980 35992 1490 36008
rect 352 35946 858 35962
rect 352 35912 858 35946
rect 352 35896 858 35912
rect 980 35850 1490 35866
rect 980 35816 1490 35850
rect 980 35800 1490 35816
rect 352 35754 858 35770
rect 352 35720 858 35754
rect 352 35704 858 35720
rect 980 35658 1490 35674
rect 980 35624 1490 35658
rect 980 35608 1490 35624
rect 352 35562 858 35578
rect 352 35528 858 35562
rect 352 35512 858 35528
rect 980 35466 1490 35482
rect 980 35432 1490 35466
rect 980 35416 1490 35432
rect 352 35370 858 35386
rect 352 35336 858 35370
rect 352 35320 858 35336
rect 980 35274 1490 35290
rect 980 35240 1490 35274
rect 980 35224 1490 35240
rect 352 35178 858 35194
rect 352 35144 858 35178
rect 352 35128 858 35144
rect 980 35082 1490 35098
rect 980 35048 1490 35082
rect 980 35032 1490 35048
rect 352 34986 858 35002
rect 352 34952 858 34986
rect 352 34936 858 34952
rect 980 34890 1490 34906
rect 980 34856 1490 34890
rect 980 34840 1490 34856
rect 352 34794 858 34810
rect 352 34760 858 34794
rect 352 34744 858 34760
rect 980 34698 1490 34714
rect 980 34664 1490 34698
rect 980 34648 1490 34664
rect 352 34602 858 34618
rect 352 34568 858 34602
rect 352 34552 858 34568
rect 980 34506 1490 34522
rect 980 34472 1490 34506
rect 980 34456 1490 34472
rect 352 34410 858 34426
rect 352 34376 858 34410
rect 352 34360 858 34376
rect 980 34314 1490 34330
rect 980 34280 1490 34314
rect 980 34264 1490 34280
rect 352 34218 858 34234
rect 352 34184 858 34218
rect 352 34168 858 34184
rect 980 34122 1490 34138
rect 980 34088 1490 34122
rect 980 34072 1490 34088
rect 352 34026 858 34042
rect 352 33992 858 34026
rect 352 33976 858 33992
rect 980 33930 1490 33946
rect 980 33896 1490 33930
rect 980 33880 1490 33896
rect 352 33834 858 33850
rect 352 33800 858 33834
rect 352 33784 858 33800
rect 980 33738 1490 33754
rect 980 33704 1490 33738
rect 980 33688 1490 33704
rect 352 33642 858 33658
rect 352 33608 858 33642
rect 352 33592 858 33608
rect 980 33546 1490 33562
rect 980 33512 1490 33546
rect 980 33496 1490 33512
rect 352 33450 858 33466
rect 352 33416 858 33450
rect 352 33400 858 33416
rect 980 33354 1490 33370
rect 980 33320 1490 33354
rect 980 33304 1490 33320
rect 352 33258 858 33274
rect 352 33224 858 33258
rect 352 33208 858 33224
rect 980 33162 1490 33178
rect 980 33128 1490 33162
rect 980 33112 1490 33128
rect 352 33066 858 33082
rect 352 33032 858 33066
rect 352 33016 858 33032
rect 980 32970 1490 32986
rect 980 32936 1490 32970
rect 980 32920 1490 32936
rect 352 32874 858 32890
rect 352 32840 858 32874
rect 352 32824 858 32840
rect 980 32778 1490 32794
rect 980 32744 1490 32778
rect 980 32728 1490 32744
rect 352 32682 858 32698
rect 352 32648 858 32682
rect 352 32632 858 32648
rect 980 32586 1490 32602
rect 980 32552 1490 32586
rect 980 32536 1490 32552
rect 352 32490 858 32506
rect 352 32456 858 32490
rect 352 32440 858 32456
rect 980 32394 1490 32410
rect 980 32360 1490 32394
rect 980 32344 1490 32360
rect 352 32298 858 32314
rect 352 32264 858 32298
rect 352 32248 858 32264
rect 980 32202 1490 32218
rect 980 32168 1490 32202
rect 980 32152 1490 32168
rect 352 32106 858 32122
rect 352 32072 858 32106
rect 352 32056 858 32072
rect 980 32010 1490 32026
rect 980 31976 1490 32010
rect 980 31960 1490 31976
rect 352 31914 858 31930
rect 352 31880 858 31914
rect 352 31864 858 31880
rect 980 31818 1490 31834
rect 980 31784 1490 31818
rect 980 31768 1490 31784
rect 352 31722 858 31738
rect 352 31688 858 31722
rect 352 31672 858 31688
rect 980 31626 1490 31642
rect 980 31592 1490 31626
rect 980 31576 1490 31592
rect 352 31530 858 31546
rect 352 31496 858 31530
rect 352 31480 858 31496
rect 980 31434 1490 31450
rect 980 31400 1490 31434
rect 980 31384 1490 31400
rect 352 31338 858 31354
rect 352 31304 858 31338
rect 352 31288 858 31304
rect 980 31242 1490 31258
rect 980 31208 1490 31242
rect 980 31192 1490 31208
rect 352 31146 858 31162
rect 352 31112 858 31146
rect 352 31096 858 31112
rect 980 31050 1490 31066
rect 980 31016 1490 31050
rect 980 31000 1490 31016
rect 352 30954 858 30970
rect 352 30920 858 30954
rect 352 30904 858 30920
rect 980 30858 1490 30874
rect 980 30824 1490 30858
rect 980 30808 1490 30824
rect 352 30762 858 30778
rect 352 30728 858 30762
rect 352 30712 858 30728
rect 980 30666 1490 30682
rect 980 30632 1490 30666
rect 980 30616 1490 30632
rect 352 30570 858 30586
rect 352 30536 858 30570
rect 352 30520 858 30536
rect 980 30474 1490 30490
rect 980 30440 1490 30474
rect 980 30424 1490 30440
rect 352 30378 858 30394
rect 352 30344 858 30378
rect 352 30328 858 30344
rect 980 30282 1490 30298
rect 980 30248 1490 30282
rect 980 30232 1490 30248
rect 352 30186 858 30202
rect 352 30152 858 30186
rect 352 30136 858 30152
rect 980 30090 1490 30106
rect 980 30056 1490 30090
rect 980 30040 1490 30056
rect 352 29994 858 30010
rect 352 29960 858 29994
rect 352 29944 858 29960
rect 980 29898 1490 29914
rect 980 29864 1490 29898
rect 980 29848 1490 29864
rect 352 29802 858 29818
rect 352 29768 858 29802
rect 352 29752 858 29768
rect 980 29706 1490 29722
rect 980 29672 1490 29706
rect 980 29656 1490 29672
rect 352 29610 858 29626
rect 352 29576 858 29610
rect 352 29560 858 29576
rect 980 29514 1490 29530
rect 980 29480 1490 29514
rect 980 29464 1490 29480
rect 352 29418 858 29434
rect 352 29384 858 29418
rect 352 29368 858 29384
rect 980 29322 1490 29338
rect 980 29288 1490 29322
rect 980 29272 1490 29288
rect 352 29226 858 29242
rect 352 29192 858 29226
rect 352 29176 858 29192
rect 980 29130 1490 29146
rect 980 29096 1490 29130
rect 980 29080 1490 29096
rect 352 29034 858 29050
rect 352 29000 858 29034
rect 352 28984 858 29000
rect 980 28938 1490 28954
rect 980 28904 1490 28938
rect 980 28888 1490 28904
rect 352 28842 858 28858
rect 352 28808 858 28842
rect 352 28792 858 28808
rect 980 28746 1490 28762
rect 980 28712 1490 28746
rect 980 28696 1490 28712
rect 352 28650 858 28666
rect 352 28616 858 28650
rect 352 28600 858 28616
rect 980 28554 1490 28570
rect 980 28520 1490 28554
rect 980 28504 1490 28520
rect 352 28458 858 28474
rect 352 28424 858 28458
rect 352 28408 858 28424
rect 980 28362 1490 28378
rect 980 28328 1490 28362
rect 980 28312 1490 28328
rect 352 28266 858 28282
rect 352 28232 858 28266
rect 352 28216 858 28232
rect 980 28170 1490 28186
rect 980 28136 1490 28170
rect 980 28120 1490 28136
rect 352 28074 858 28090
rect 352 28040 858 28074
rect 352 28024 858 28040
rect 980 27978 1490 27994
rect 980 27944 1490 27978
rect 980 27928 1490 27944
rect 352 27882 858 27898
rect 352 27848 858 27882
rect 352 27832 858 27848
rect 980 27786 1490 27802
rect 980 27752 1490 27786
rect 980 27736 1490 27752
rect 352 27690 858 27706
rect 352 27656 858 27690
rect 352 27640 858 27656
rect 980 27594 1490 27610
rect 980 27560 1490 27594
rect 980 27544 1490 27560
rect 352 27498 858 27514
rect 352 27464 858 27498
rect 352 27448 858 27464
rect 980 27402 1490 27418
rect 980 27368 1490 27402
rect 980 27352 1490 27368
rect 352 27306 858 27322
rect 352 27272 858 27306
rect 352 27256 858 27272
rect 980 27210 1490 27226
rect 980 27176 1490 27210
rect 980 27160 1490 27176
rect 352 27114 858 27130
rect 352 27080 858 27114
rect 352 27064 858 27080
rect 980 27018 1490 27034
rect 980 26984 1490 27018
rect 980 26968 1490 26984
rect 352 26922 858 26938
rect 352 26888 858 26922
rect 352 26872 858 26888
rect 980 26826 1490 26842
rect 980 26792 1490 26826
rect 980 26776 1490 26792
rect 352 26730 858 26746
rect 352 26696 858 26730
rect 352 26680 858 26696
rect 980 26634 1490 26650
rect 980 26600 1490 26634
rect 980 26584 1490 26600
rect 352 26538 858 26554
rect 352 26504 858 26538
rect 352 26488 858 26504
rect 980 26442 1490 26458
rect 980 26408 1490 26442
rect 980 26392 1490 26408
rect 352 26346 858 26362
rect 352 26312 858 26346
rect 352 26296 858 26312
rect 980 26250 1490 26266
rect 980 26216 1490 26250
rect 980 26200 1490 26216
rect 352 26154 858 26170
rect 352 26120 858 26154
rect 352 26104 858 26120
rect 980 26058 1490 26074
rect 980 26024 1490 26058
rect 980 26008 1490 26024
rect 352 25962 858 25978
rect 352 25928 858 25962
rect 352 25912 858 25928
rect 980 25866 1490 25882
rect 980 25832 1490 25866
rect 980 25816 1490 25832
rect 352 25770 858 25786
rect 352 25736 858 25770
rect 352 25720 858 25736
rect 980 25674 1490 25690
rect 980 25640 1490 25674
rect 980 25624 1490 25640
rect 352 25578 858 25594
rect 352 25544 858 25578
rect 352 25528 858 25544
rect 980 25482 1490 25498
rect 980 25448 1490 25482
rect 980 25432 1490 25448
rect 352 25386 858 25402
rect 352 25352 858 25386
rect 352 25336 858 25352
rect 980 25290 1490 25306
rect 980 25256 1490 25290
rect 980 25240 1490 25256
rect 352 25194 858 25210
rect 352 25160 858 25194
rect 352 25144 858 25160
rect 980 25098 1490 25114
rect 980 25064 1490 25098
rect 980 25048 1490 25064
rect 352 25002 858 25018
rect 352 24968 858 25002
rect 352 24952 858 24968
rect 980 24906 1490 24922
rect 980 24872 1490 24906
rect 980 24856 1490 24872
rect 352 24810 858 24826
rect 352 24776 858 24810
rect 352 24760 858 24776
rect 980 24714 1490 24730
rect 980 24680 1490 24714
rect 980 24664 1490 24680
rect 352 24618 858 24634
rect 352 24584 858 24618
rect 352 24568 858 24584
rect 980 24522 1490 24538
rect 980 24488 1490 24522
rect 980 24472 1490 24488
rect 352 24426 858 24442
rect 352 24392 858 24426
rect 352 24376 858 24392
rect 980 24330 1490 24346
rect 980 24296 1490 24330
rect 980 24280 1490 24296
rect 352 24234 858 24250
rect 352 24200 858 24234
rect 352 24184 858 24200
rect 980 24138 1490 24154
rect 980 24104 1490 24138
rect 980 24088 1490 24104
rect 352 24042 858 24058
rect 352 24008 858 24042
rect 352 23992 858 24008
rect 980 23946 1490 23962
rect 980 23912 1490 23946
rect 980 23896 1490 23912
rect 352 23850 858 23866
rect 352 23816 858 23850
rect 352 23800 858 23816
rect 980 23754 1490 23770
rect 980 23720 1490 23754
rect 980 23704 1490 23720
rect 352 23658 858 23674
rect 352 23624 858 23658
rect 352 23608 858 23624
rect 980 23562 1490 23578
rect 980 23528 1490 23562
rect 980 23512 1490 23528
rect 352 23466 858 23482
rect 352 23432 858 23466
rect 352 23416 858 23432
rect 980 23370 1490 23386
rect 980 23336 1490 23370
rect 980 23320 1490 23336
rect 352 23274 858 23290
rect 352 23240 858 23274
rect 352 23224 858 23240
rect 980 23178 1490 23194
rect 980 23144 1490 23178
rect 980 23128 1490 23144
rect 352 23082 858 23098
rect 352 23048 858 23082
rect 352 23032 858 23048
rect 340 21986 870 22768
rect 352 21704 858 21720
rect 352 21670 858 21704
rect 352 21654 858 21670
rect 980 21608 1490 21624
rect 980 21574 1490 21608
rect 980 21558 1490 21574
rect 352 21512 858 21528
rect 352 21478 858 21512
rect 352 21462 858 21478
rect 980 21416 1490 21432
rect 980 21382 1490 21416
rect 980 21366 1490 21382
rect 352 21320 858 21336
rect 352 21286 858 21320
rect 352 21270 858 21286
rect 980 21224 1490 21240
rect 980 21190 1490 21224
rect 980 21174 1490 21190
rect 352 21128 858 21144
rect 352 21094 858 21128
rect 352 21078 858 21094
rect 980 21032 1490 21048
rect 980 20998 1490 21032
rect 980 20982 1490 20998
rect 352 20936 858 20952
rect 352 20902 858 20936
rect 352 20886 858 20902
rect 980 20840 1490 20856
rect 980 20806 1490 20840
rect 980 20790 1490 20806
rect 352 20744 858 20760
rect 352 20710 858 20744
rect 352 20694 858 20710
rect 980 20648 1490 20664
rect 980 20614 1490 20648
rect 980 20598 1490 20614
rect 352 20552 858 20568
rect 352 20518 858 20552
rect 352 20502 858 20518
rect 980 20456 1490 20472
rect 980 20422 1490 20456
rect 980 20406 1490 20422
rect 352 20360 858 20376
rect 352 20326 858 20360
rect 352 20310 858 20326
rect 980 20264 1490 20280
rect 980 20230 1490 20264
rect 980 20214 1490 20230
rect 352 20168 858 20184
rect 352 20134 858 20168
rect 352 20118 858 20134
rect 980 20072 1490 20088
rect 980 20038 1490 20072
rect 980 20022 1490 20038
rect 352 19976 858 19992
rect 352 19942 858 19976
rect 352 19926 858 19942
rect 980 19880 1490 19896
rect 980 19846 1490 19880
rect 980 19830 1490 19846
rect 352 19784 858 19800
rect 352 19750 858 19784
rect 352 19734 858 19750
rect 980 19688 1490 19704
rect 980 19654 1490 19688
rect 980 19638 1490 19654
rect 352 19592 858 19608
rect 352 19558 858 19592
rect 352 19542 858 19558
rect 980 19496 1490 19512
rect 980 19462 1490 19496
rect 980 19446 1490 19462
rect 352 19400 858 19416
rect 352 19366 858 19400
rect 352 19350 858 19366
rect 980 19304 1490 19320
rect 980 19270 1490 19304
rect 980 19254 1490 19270
rect 352 19208 858 19224
rect 352 19174 858 19208
rect 352 19158 858 19174
rect 980 19112 1490 19128
rect 980 19078 1490 19112
rect 980 19062 1490 19078
rect 352 19016 858 19032
rect 352 18982 858 19016
rect 352 18966 858 18982
rect 980 18920 1490 18936
rect 980 18886 1490 18920
rect 980 18870 1490 18886
rect 352 18824 858 18840
rect 352 18790 858 18824
rect 352 18774 858 18790
rect 980 18728 1490 18744
rect 980 18694 1490 18728
rect 980 18678 1490 18694
rect 352 18632 858 18648
rect 352 18598 858 18632
rect 352 18582 858 18598
rect 980 18536 1490 18552
rect 980 18502 1490 18536
rect 980 18486 1490 18502
rect 352 18440 858 18456
rect 352 18406 858 18440
rect 352 18390 858 18406
rect 980 18344 1490 18360
rect 980 18310 1490 18344
rect 980 18294 1490 18310
rect 352 18248 858 18264
rect 352 18214 858 18248
rect 352 18198 858 18214
rect 980 18152 1490 18168
rect 980 18118 1490 18152
rect 980 18102 1490 18118
rect 352 18056 858 18072
rect 352 18022 858 18056
rect 352 18006 858 18022
rect 980 17960 1490 17976
rect 980 17926 1490 17960
rect 980 17910 1490 17926
rect 352 17864 858 17880
rect 352 17830 858 17864
rect 352 17814 858 17830
rect 980 17768 1490 17784
rect 980 17734 1490 17768
rect 980 17718 1490 17734
rect 352 17672 858 17688
rect 352 17638 858 17672
rect 352 17622 858 17638
rect 980 17576 1490 17592
rect 980 17542 1490 17576
rect 980 17526 1490 17542
rect 352 17480 858 17496
rect 352 17446 858 17480
rect 352 17430 858 17446
rect 980 17384 1490 17400
rect 980 17350 1490 17384
rect 980 17334 1490 17350
rect 352 17288 858 17304
rect 352 17254 858 17288
rect 352 17238 858 17254
rect 980 17192 1490 17208
rect 980 17158 1490 17192
rect 980 17142 1490 17158
rect 352 17096 858 17112
rect 352 17062 858 17096
rect 352 17046 858 17062
rect 980 17000 1490 17016
rect 980 16966 1490 17000
rect 980 16950 1490 16966
rect 352 16904 858 16920
rect 352 16870 858 16904
rect 352 16854 858 16870
rect 980 16808 1490 16824
rect 980 16774 1490 16808
rect 980 16758 1490 16774
rect 352 16712 858 16728
rect 352 16678 858 16712
rect 352 16662 858 16678
rect 980 16616 1490 16632
rect 980 16582 1490 16616
rect 980 16566 1490 16582
rect 352 16520 858 16536
rect 352 16486 858 16520
rect 352 16470 858 16486
rect 980 16424 1490 16440
rect 980 16390 1490 16424
rect 980 16374 1490 16390
rect 352 16328 858 16344
rect 352 16294 858 16328
rect 352 16278 858 16294
rect 980 16232 1490 16248
rect 980 16198 1490 16232
rect 980 16182 1490 16198
rect 352 16136 858 16152
rect 352 16102 858 16136
rect 352 16086 858 16102
rect 980 16040 1490 16056
rect 980 16006 1490 16040
rect 980 15990 1490 16006
rect 352 15944 858 15960
rect 352 15910 858 15944
rect 352 15894 858 15910
rect 980 15848 1490 15864
rect 980 15814 1490 15848
rect 980 15798 1490 15814
rect 352 15752 858 15768
rect 352 15718 858 15752
rect 352 15702 858 15718
rect 980 15656 1490 15672
rect 980 15622 1490 15656
rect 980 15606 1490 15622
rect 352 15560 858 15576
rect 352 15526 858 15560
rect 352 15510 858 15526
rect 980 15464 1490 15480
rect 980 15430 1490 15464
rect 980 15414 1490 15430
rect 352 15368 858 15384
rect 352 15334 858 15368
rect 352 15318 858 15334
rect 980 15272 1490 15288
rect 980 15238 1490 15272
rect 980 15222 1490 15238
rect 352 15176 858 15192
rect 352 15142 858 15176
rect 352 15126 858 15142
rect 980 15080 1490 15096
rect 980 15046 1490 15080
rect 980 15030 1490 15046
rect 352 14984 858 15000
rect 352 14950 858 14984
rect 352 14934 858 14950
rect 980 14888 1490 14904
rect 980 14854 1490 14888
rect 980 14838 1490 14854
rect 352 14792 858 14808
rect 352 14758 858 14792
rect 352 14742 858 14758
rect 980 14696 1490 14712
rect 980 14662 1490 14696
rect 980 14646 1490 14662
rect 352 14600 858 14616
rect 352 14566 858 14600
rect 352 14550 858 14566
rect 980 14504 1490 14520
rect 980 14470 1490 14504
rect 980 14454 1490 14470
rect 352 14408 858 14424
rect 352 14374 858 14408
rect 352 14358 858 14374
rect 980 14312 1490 14328
rect 980 14278 1490 14312
rect 980 14262 1490 14278
rect 352 14216 858 14232
rect 352 14182 858 14216
rect 352 14166 858 14182
rect 980 14120 1490 14136
rect 980 14086 1490 14120
rect 980 14070 1490 14086
rect 352 14024 858 14040
rect 352 13990 858 14024
rect 352 13974 858 13990
rect 980 13928 1490 13944
rect 980 13894 1490 13928
rect 980 13878 1490 13894
rect 352 13832 858 13848
rect 352 13798 858 13832
rect 352 13782 858 13798
rect 980 13736 1490 13752
rect 980 13702 1490 13736
rect 980 13686 1490 13702
rect 352 13640 858 13656
rect 352 13606 858 13640
rect 352 13590 858 13606
rect 980 13544 1490 13560
rect 980 13510 1490 13544
rect 980 13494 1490 13510
rect 352 13448 858 13464
rect 352 13414 858 13448
rect 352 13398 858 13414
rect 980 13352 1490 13368
rect 980 13318 1490 13352
rect 980 13302 1490 13318
rect 352 13256 858 13272
rect 352 13222 858 13256
rect 352 13206 858 13222
rect 980 13160 1490 13176
rect 980 13126 1490 13160
rect 980 13110 1490 13126
rect 352 13064 858 13080
rect 352 13030 858 13064
rect 352 13014 858 13030
rect 980 12968 1490 12984
rect 980 12934 1490 12968
rect 980 12918 1490 12934
rect 352 12872 858 12888
rect 352 12838 858 12872
rect 352 12822 858 12838
rect 980 12776 1490 12792
rect 980 12742 1490 12776
rect 980 12726 1490 12742
rect 352 12680 858 12696
rect 352 12646 858 12680
rect 352 12630 858 12646
rect 980 12584 1490 12600
rect 980 12550 1490 12584
rect 980 12534 1490 12550
rect 352 12488 858 12504
rect 352 12454 858 12488
rect 352 12438 858 12454
rect 980 12392 1490 12408
rect 980 12358 1490 12392
rect 980 12342 1490 12358
rect 352 12296 858 12312
rect 352 12262 858 12296
rect 352 12246 858 12262
rect 980 12200 1490 12216
rect 980 12166 1490 12200
rect 980 12150 1490 12166
rect 352 12104 858 12120
rect 352 12070 858 12104
rect 352 12054 858 12070
rect 980 12008 1490 12024
rect 980 11974 1490 12008
rect 980 11958 1490 11974
rect 352 11912 858 11928
rect 352 11878 858 11912
rect 352 11862 858 11878
rect 980 11816 1490 11832
rect 980 11782 1490 11816
rect 980 11766 1490 11782
rect 352 11720 858 11736
rect 352 11686 858 11720
rect 352 11670 858 11686
rect 980 11624 1490 11640
rect 980 11590 1490 11624
rect 980 11574 1490 11590
rect 352 11528 858 11544
rect 352 11494 858 11528
rect 352 11478 858 11494
rect 980 11432 1490 11448
rect 980 11398 1490 11432
rect 980 11382 1490 11398
rect 352 11336 858 11352
rect 352 11302 858 11336
rect 352 11286 858 11302
rect 980 11240 1490 11256
rect 980 11206 1490 11240
rect 980 11190 1490 11206
rect 352 11144 858 11160
rect 352 11110 858 11144
rect 352 11094 858 11110
rect 980 11048 1490 11064
rect 980 11014 1490 11048
rect 980 10998 1490 11014
rect 352 10952 858 10968
rect 352 10918 858 10952
rect 352 10902 858 10918
rect 980 10856 1490 10872
rect 980 10822 1490 10856
rect 980 10806 1490 10822
rect 352 10760 858 10776
rect 352 10726 858 10760
rect 352 10710 858 10726
rect 980 10664 1490 10680
rect 980 10630 1490 10664
rect 980 10614 1490 10630
rect 352 10568 858 10584
rect 352 10534 858 10568
rect 352 10518 858 10534
rect 980 10472 1490 10488
rect 980 10438 1490 10472
rect 980 10422 1490 10438
rect 352 10376 858 10392
rect 352 10342 858 10376
rect 352 10326 858 10342
rect 980 10280 1490 10296
rect 980 10246 1490 10280
rect 980 10230 1490 10246
rect 352 10184 858 10200
rect 352 10150 858 10184
rect 352 10134 858 10150
rect 980 10088 1490 10104
rect 980 10054 1490 10088
rect 980 10038 1490 10054
rect 352 9992 858 10008
rect 352 9958 858 9992
rect 352 9942 858 9958
rect 980 9896 1490 9912
rect 980 9862 1490 9896
rect 980 9846 1490 9862
rect 352 9800 858 9816
rect 352 9766 858 9800
rect 352 9750 858 9766
rect 980 9704 1490 9720
rect 980 9670 1490 9704
rect 980 9654 1490 9670
rect 352 9608 858 9624
rect 352 9574 858 9608
rect 352 9558 858 9574
rect 980 9512 1490 9528
rect 980 9478 1490 9512
rect 980 9462 1490 9478
rect 352 9416 858 9432
rect 352 9382 858 9416
rect 352 9366 858 9382
rect 980 9320 1490 9336
rect 980 9286 1490 9320
rect 980 9270 1490 9286
rect 352 9224 858 9240
rect 352 9190 858 9224
rect 352 9174 858 9190
rect 980 9128 1490 9144
rect 980 9094 1490 9128
rect 980 9078 1490 9094
rect 352 9032 858 9048
rect 352 8998 858 9032
rect 352 8982 858 8998
rect 980 8936 1490 8952
rect 980 8902 1490 8936
rect 980 8886 1490 8902
rect 352 8840 858 8856
rect 352 8806 858 8840
rect 352 8790 858 8806
rect 980 8744 1490 8760
rect 980 8710 1490 8744
rect 980 8694 1490 8710
rect 352 8648 858 8664
rect 352 8614 858 8648
rect 352 8598 858 8614
rect 980 8552 1490 8568
rect 980 8518 1490 8552
rect 980 8502 1490 8518
rect 352 8456 858 8472
rect 352 8422 858 8456
rect 352 8406 858 8422
rect 980 8360 1490 8376
rect 980 8326 1490 8360
rect 980 8310 1490 8326
rect 352 8264 858 8280
rect 352 8230 858 8264
rect 352 8214 858 8230
rect 980 8168 1490 8184
rect 980 8134 1490 8168
rect 980 8118 1490 8134
rect 352 8072 858 8088
rect 352 8038 858 8072
rect 352 8022 858 8038
rect 980 7976 1490 7992
rect 980 7942 1490 7976
rect 980 7926 1490 7942
rect 352 7880 858 7896
rect 352 7846 858 7880
rect 352 7830 858 7846
rect 980 7784 1490 7800
rect 980 7750 1490 7784
rect 980 7734 1490 7750
rect 352 7688 858 7704
rect 352 7654 858 7688
rect 352 7638 858 7654
rect 980 7592 1490 7608
rect 980 7558 1490 7592
rect 980 7542 1490 7558
rect 352 7496 858 7512
rect 352 7462 858 7496
rect 352 7446 858 7462
rect 980 7400 1490 7416
rect 980 7366 1490 7400
rect 980 7350 1490 7366
rect 352 7304 858 7320
rect 352 7270 858 7304
rect 352 7254 858 7270
rect 980 7208 1490 7224
rect 980 7174 1490 7208
rect 980 7158 1490 7174
rect 352 7112 858 7128
rect 352 7078 858 7112
rect 352 7062 858 7078
rect 980 7016 1490 7032
rect 980 6982 1490 7016
rect 980 6966 1490 6982
rect 352 6920 858 6936
rect 352 6886 858 6920
rect 352 6870 858 6886
rect 980 6824 1490 6840
rect 980 6790 1490 6824
rect 980 6774 1490 6790
rect 352 6728 858 6744
rect 352 6694 858 6728
rect 352 6678 858 6694
rect 980 6632 1490 6648
rect 980 6598 1490 6632
rect 980 6582 1490 6598
rect 352 6536 858 6552
rect 352 6502 858 6536
rect 352 6486 858 6502
rect 980 6440 1490 6456
rect 980 6406 1490 6440
rect 980 6390 1490 6406
rect 352 6344 858 6360
rect 352 6310 858 6344
rect 352 6294 858 6310
rect 980 6248 1490 6264
rect 980 6214 1490 6248
rect 980 6198 1490 6214
rect 352 6152 858 6168
rect 352 6118 858 6152
rect 352 6102 858 6118
rect 980 6056 1490 6072
rect 980 6022 1490 6056
rect 980 6006 1490 6022
rect 352 5960 858 5976
rect 352 5926 858 5960
rect 352 5910 858 5926
rect 980 5864 1490 5880
rect 980 5830 1490 5864
rect 980 5814 1490 5830
rect 352 5768 858 5784
rect 352 5734 858 5768
rect 352 5718 858 5734
rect 980 5672 1490 5688
rect 980 5638 1490 5672
rect 980 5622 1490 5638
rect 352 5576 858 5592
rect 352 5542 858 5576
rect 352 5526 858 5542
rect 980 5480 1490 5496
rect 980 5446 1490 5480
rect 980 5430 1490 5446
rect 352 5384 858 5400
rect 352 5350 858 5384
rect 352 5334 858 5350
rect 980 5288 1490 5304
rect 980 5254 1490 5288
rect 980 5238 1490 5254
rect 352 5192 858 5208
rect 352 5158 858 5192
rect 352 5142 858 5158
rect 980 5096 1490 5112
rect 980 5062 1490 5096
rect 980 5046 1490 5062
rect 352 5000 858 5016
rect 352 4966 858 5000
rect 352 4950 858 4966
rect 980 4904 1490 4920
rect 980 4870 1490 4904
rect 980 4854 1490 4870
rect 352 4808 858 4824
rect 352 4774 858 4808
rect 352 4758 858 4774
rect 980 4712 1490 4728
rect 980 4678 1490 4712
rect 980 4662 1490 4678
rect 352 4616 858 4632
rect 352 4582 858 4616
rect 352 4566 858 4582
rect 980 4520 1490 4536
rect 980 4486 1490 4520
rect 980 4470 1490 4486
rect 352 4424 858 4440
rect 352 4390 858 4424
rect 352 4374 858 4390
rect 980 4328 1490 4344
rect 980 4294 1490 4328
rect 980 4278 1490 4294
rect 352 4232 858 4248
rect 352 4198 858 4232
rect 352 4182 858 4198
rect 980 4136 1490 4152
rect 980 4102 1490 4136
rect 980 4086 1490 4102
rect 352 4040 858 4056
rect 352 4006 858 4040
rect 352 3990 858 4006
rect 980 3944 1490 3960
rect 980 3910 1490 3944
rect 980 3894 1490 3910
rect 352 3848 858 3864
rect 352 3814 858 3848
rect 352 3798 858 3814
rect 980 3752 1490 3768
rect 980 3718 1490 3752
rect 980 3702 1490 3718
rect 352 3656 858 3672
rect 352 3622 858 3656
rect 352 3606 858 3622
rect 980 3560 1490 3576
rect 980 3526 1490 3560
rect 980 3510 1490 3526
rect 352 3464 858 3480
rect 352 3430 858 3464
rect 352 3414 858 3430
rect 980 3368 1490 3384
rect 980 3334 1490 3368
rect 980 3318 1490 3334
rect 352 3272 858 3288
rect 352 3238 858 3272
rect 352 3222 858 3238
rect 980 3176 1490 3192
rect 980 3142 1490 3176
rect 980 3126 1490 3142
rect 352 3080 858 3096
rect 352 3046 858 3080
rect 352 3030 858 3046
rect 980 2984 1490 3000
rect 980 2950 1490 2984
rect 980 2934 1490 2950
rect 352 2888 858 2904
rect 352 2854 858 2888
rect 352 2838 858 2854
rect 980 2792 1490 2808
rect 980 2758 1490 2792
rect 980 2742 1490 2758
rect 352 2696 858 2712
rect 352 2662 858 2696
rect 352 2646 858 2662
rect 980 2600 1490 2616
rect 980 2566 1490 2600
rect 980 2550 1490 2566
rect 352 2504 858 2520
rect 352 2470 858 2504
rect 352 2454 858 2470
rect 980 2408 1490 2424
rect 980 2374 1490 2408
rect 980 2358 1490 2374
rect 352 2312 858 2328
rect 352 2278 858 2312
rect 352 2262 858 2278
rect 980 2216 1490 2232
rect 980 2182 1490 2216
rect 980 2166 1490 2182
rect 352 2120 858 2136
rect 352 2086 858 2120
rect 352 2070 858 2086
rect 980 2024 1490 2040
rect 980 1990 1490 2024
rect 980 1974 1490 1990
rect 352 1928 858 1944
rect 352 1894 858 1928
rect 352 1878 858 1894
rect 980 1832 1490 1848
rect 980 1798 1490 1832
rect 980 1782 1490 1798
rect 352 1736 858 1752
rect 352 1702 858 1736
rect 352 1686 858 1702
rect 980 1640 1490 1656
rect 980 1606 1490 1640
rect 980 1590 1490 1606
rect 352 1544 858 1560
rect 352 1510 858 1544
rect 352 1494 858 1510
rect 980 1448 1490 1464
rect 980 1414 1490 1448
rect 980 1398 1490 1414
rect 352 1352 858 1368
rect 352 1318 858 1352
rect 352 1302 858 1318
rect 980 1256 1490 1272
rect 980 1222 1490 1256
rect 980 1206 1490 1222
rect 352 1160 858 1176
rect 352 1126 858 1160
rect 352 1110 858 1126
rect 980 1064 1490 1080
rect 980 1030 1490 1064
rect 980 1014 1490 1030
rect 352 968 858 984
rect 352 934 858 968
rect 352 918 858 934
rect 980 872 1490 888
rect 980 838 1490 872
rect 980 822 1490 838
rect 352 776 858 792
rect 352 742 858 776
rect 352 726 858 742
rect 980 680 1490 696
rect 980 646 1490 680
rect 980 630 1490 646
rect 352 584 858 600
rect 352 550 858 584
rect 352 534 858 550
<< metal2 >>
rect 132 45136 1706 45146
rect 132 45052 1706 45062
rect 342 44218 868 44228
rect 342 44152 352 44218
rect 858 44152 868 44218
rect 342 44142 868 44152
rect 970 44122 1500 44132
rect 970 44056 980 44122
rect 1490 44056 1500 44122
rect 970 44046 1500 44056
rect 342 44026 868 44036
rect 342 43960 352 44026
rect 858 43960 868 44026
rect 342 43950 868 43960
rect 970 43930 1500 43940
rect 970 43864 980 43930
rect 1490 43864 1500 43930
rect 970 43854 1500 43864
rect 342 43834 868 43844
rect 342 43768 352 43834
rect 858 43768 868 43834
rect 342 43758 868 43768
rect 970 43738 1500 43748
rect 970 43672 980 43738
rect 1490 43672 1500 43738
rect 970 43662 1500 43672
rect 342 43642 868 43652
rect 342 43576 352 43642
rect 858 43576 868 43642
rect 342 43566 868 43576
rect 970 43546 1500 43556
rect 970 43480 980 43546
rect 1490 43480 1500 43546
rect 970 43470 1500 43480
rect 342 43450 868 43460
rect 342 43384 352 43450
rect 858 43384 868 43450
rect 342 43374 868 43384
rect 970 43354 1500 43364
rect 970 43288 980 43354
rect 1490 43288 1500 43354
rect 970 43278 1500 43288
rect 342 43258 868 43268
rect 342 43192 352 43258
rect 858 43192 868 43258
rect 342 43182 868 43192
rect 970 43162 1500 43172
rect 970 43096 980 43162
rect 1490 43096 1500 43162
rect 970 43086 1500 43096
rect 342 43066 868 43076
rect 342 43000 352 43066
rect 858 43000 868 43066
rect 342 42990 868 43000
rect 970 42970 1500 42980
rect 970 42904 980 42970
rect 1490 42904 1500 42970
rect 970 42894 1500 42904
rect 342 42874 868 42884
rect 342 42808 352 42874
rect 858 42808 868 42874
rect 342 42798 868 42808
rect 970 42778 1500 42788
rect 970 42712 980 42778
rect 1490 42712 1500 42778
rect 970 42702 1500 42712
rect 342 42682 868 42692
rect 342 42616 352 42682
rect 858 42616 868 42682
rect 342 42606 868 42616
rect 970 42586 1500 42596
rect 970 42520 980 42586
rect 1490 42520 1500 42586
rect 970 42510 1500 42520
rect 342 42490 868 42500
rect 342 42424 352 42490
rect 858 42424 868 42490
rect 342 42414 868 42424
rect 970 42394 1500 42404
rect 970 42328 980 42394
rect 1490 42328 1500 42394
rect 970 42318 1500 42328
rect 342 42298 868 42308
rect 342 42232 352 42298
rect 858 42232 868 42298
rect 342 42222 868 42232
rect 970 42202 1500 42212
rect 970 42136 980 42202
rect 1490 42136 1500 42202
rect 970 42126 1500 42136
rect 342 42106 868 42116
rect 342 42040 352 42106
rect 858 42040 868 42106
rect 342 42030 868 42040
rect 970 42010 1500 42020
rect 970 41944 980 42010
rect 1490 41944 1500 42010
rect 970 41934 1500 41944
rect 342 41914 868 41924
rect 342 41848 352 41914
rect 858 41848 868 41914
rect 342 41838 868 41848
rect 970 41818 1500 41828
rect 970 41752 980 41818
rect 1490 41752 1500 41818
rect 970 41742 1500 41752
rect 342 41722 868 41732
rect 342 41656 352 41722
rect 858 41656 868 41722
rect 342 41646 868 41656
rect 970 41626 1500 41636
rect 970 41560 980 41626
rect 1490 41560 1500 41626
rect 970 41550 1500 41560
rect 342 41530 868 41540
rect 342 41464 352 41530
rect 858 41464 868 41530
rect 342 41454 868 41464
rect 970 41434 1500 41444
rect 970 41368 980 41434
rect 1490 41368 1500 41434
rect 970 41358 1500 41368
rect 342 41338 868 41348
rect 342 41272 352 41338
rect 858 41272 868 41338
rect 342 41262 868 41272
rect 970 41242 1500 41252
rect 970 41176 980 41242
rect 1490 41176 1500 41242
rect 970 41166 1500 41176
rect 342 41146 868 41156
rect 342 41080 352 41146
rect 858 41080 868 41146
rect 342 41070 868 41080
rect 970 41050 1500 41060
rect 970 40984 980 41050
rect 1490 40984 1500 41050
rect 970 40974 1500 40984
rect 342 40954 868 40964
rect 342 40888 352 40954
rect 858 40888 868 40954
rect 342 40878 868 40888
rect 970 40858 1500 40868
rect 970 40792 980 40858
rect 1490 40792 1500 40858
rect 970 40782 1500 40792
rect 342 40762 868 40772
rect 342 40696 352 40762
rect 858 40696 868 40762
rect 342 40686 868 40696
rect 970 40666 1500 40676
rect 970 40600 980 40666
rect 1490 40600 1500 40666
rect 970 40590 1500 40600
rect 342 40570 868 40580
rect 342 40504 352 40570
rect 858 40504 868 40570
rect 342 40494 868 40504
rect 970 40474 1500 40484
rect 970 40408 980 40474
rect 1490 40408 1500 40474
rect 970 40398 1500 40408
rect 342 40378 868 40388
rect 342 40312 352 40378
rect 858 40312 868 40378
rect 342 40302 868 40312
rect 970 40282 1500 40292
rect 970 40216 980 40282
rect 1490 40216 1500 40282
rect 970 40206 1500 40216
rect 342 40186 868 40196
rect 342 40120 352 40186
rect 858 40120 868 40186
rect 342 40110 868 40120
rect 970 40090 1500 40100
rect 970 40024 980 40090
rect 1490 40024 1500 40090
rect 970 40014 1500 40024
rect 342 39994 868 40004
rect 342 39928 352 39994
rect 858 39928 868 39994
rect 342 39918 868 39928
rect 970 39898 1500 39908
rect 970 39832 980 39898
rect 1490 39832 1500 39898
rect 970 39822 1500 39832
rect 342 39802 868 39812
rect 342 39736 352 39802
rect 858 39736 868 39802
rect 342 39726 868 39736
rect 970 39706 1500 39716
rect 970 39640 980 39706
rect 1490 39640 1500 39706
rect 970 39630 1500 39640
rect 342 39610 868 39620
rect 342 39544 352 39610
rect 858 39544 868 39610
rect 342 39534 868 39544
rect 970 39514 1500 39524
rect 970 39448 980 39514
rect 1490 39448 1500 39514
rect 970 39438 1500 39448
rect 342 39418 868 39428
rect 342 39352 352 39418
rect 858 39352 868 39418
rect 342 39342 868 39352
rect 970 39322 1500 39332
rect 970 39256 980 39322
rect 1490 39256 1500 39322
rect 970 39246 1500 39256
rect 342 39226 868 39236
rect 342 39160 352 39226
rect 858 39160 868 39226
rect 342 39150 868 39160
rect 970 39130 1500 39140
rect 970 39064 980 39130
rect 1490 39064 1500 39130
rect 970 39054 1500 39064
rect 342 39034 868 39044
rect 342 38968 352 39034
rect 858 38968 868 39034
rect 342 38958 868 38968
rect 970 38938 1500 38948
rect 970 38872 980 38938
rect 1490 38872 1500 38938
rect 970 38862 1500 38872
rect 342 38842 868 38852
rect 342 38776 352 38842
rect 858 38776 868 38842
rect 342 38766 868 38776
rect 970 38746 1500 38756
rect 970 38680 980 38746
rect 1490 38680 1500 38746
rect 970 38670 1500 38680
rect 342 38650 868 38660
rect 342 38584 352 38650
rect 858 38584 868 38650
rect 342 38574 868 38584
rect 970 38554 1500 38564
rect 970 38488 980 38554
rect 1490 38488 1500 38554
rect 970 38478 1500 38488
rect 342 38458 868 38468
rect 342 38392 352 38458
rect 858 38392 868 38458
rect 342 38382 868 38392
rect 970 38362 1500 38372
rect 970 38296 980 38362
rect 1490 38296 1500 38362
rect 970 38286 1500 38296
rect 342 38266 868 38276
rect 342 38200 352 38266
rect 858 38200 868 38266
rect 342 38190 868 38200
rect 970 38170 1500 38180
rect 970 38104 980 38170
rect 1490 38104 1500 38170
rect 970 38094 1500 38104
rect 342 38074 868 38084
rect 342 38008 352 38074
rect 858 38008 868 38074
rect 342 37998 868 38008
rect 970 37978 1500 37988
rect 970 37912 980 37978
rect 1490 37912 1500 37978
rect 970 37902 1500 37912
rect 342 37882 868 37892
rect 342 37816 352 37882
rect 858 37816 868 37882
rect 342 37806 868 37816
rect 970 37786 1500 37796
rect 970 37720 980 37786
rect 1490 37720 1500 37786
rect 970 37710 1500 37720
rect 342 37690 868 37700
rect 342 37624 352 37690
rect 858 37624 868 37690
rect 342 37614 868 37624
rect 970 37594 1500 37604
rect 970 37528 980 37594
rect 1490 37528 1500 37594
rect 970 37518 1500 37528
rect 342 37498 868 37508
rect 342 37432 352 37498
rect 858 37432 868 37498
rect 342 37422 868 37432
rect 970 37402 1500 37412
rect 970 37336 980 37402
rect 1490 37336 1500 37402
rect 970 37326 1500 37336
rect 342 37306 868 37316
rect 342 37240 352 37306
rect 858 37240 868 37306
rect 342 37230 868 37240
rect 970 37210 1500 37220
rect 970 37144 980 37210
rect 1490 37144 1500 37210
rect 970 37134 1500 37144
rect 342 37114 868 37124
rect 342 37048 352 37114
rect 858 37048 868 37114
rect 342 37038 868 37048
rect 970 37018 1500 37028
rect 970 36952 980 37018
rect 1490 36952 1500 37018
rect 970 36942 1500 36952
rect 342 36922 868 36932
rect 342 36856 352 36922
rect 858 36856 868 36922
rect 342 36846 868 36856
rect 970 36826 1500 36836
rect 970 36760 980 36826
rect 1490 36760 1500 36826
rect 970 36750 1500 36760
rect 342 36730 868 36740
rect 342 36664 352 36730
rect 858 36664 868 36730
rect 342 36654 868 36664
rect 970 36634 1500 36644
rect 970 36568 980 36634
rect 1490 36568 1500 36634
rect 970 36558 1500 36568
rect 342 36538 868 36548
rect 342 36472 352 36538
rect 858 36472 868 36538
rect 342 36462 868 36472
rect 970 36442 1500 36452
rect 970 36376 980 36442
rect 1490 36376 1500 36442
rect 970 36366 1500 36376
rect 342 36346 868 36356
rect 342 36280 352 36346
rect 858 36280 868 36346
rect 342 36270 868 36280
rect 970 36250 1500 36260
rect 970 36184 980 36250
rect 1490 36184 1500 36250
rect 970 36174 1500 36184
rect 342 36154 868 36164
rect 342 36088 352 36154
rect 858 36088 868 36154
rect 342 36078 868 36088
rect 970 36058 1500 36068
rect 970 35992 980 36058
rect 1490 35992 1500 36058
rect 970 35982 1500 35992
rect 342 35962 868 35972
rect 342 35896 352 35962
rect 858 35896 868 35962
rect 342 35886 868 35896
rect 970 35866 1500 35876
rect 970 35800 980 35866
rect 1490 35800 1500 35866
rect 970 35790 1500 35800
rect 342 35770 868 35780
rect 342 35704 352 35770
rect 858 35704 868 35770
rect 342 35694 868 35704
rect 970 35674 1500 35684
rect 970 35608 980 35674
rect 1490 35608 1500 35674
rect 970 35598 1500 35608
rect 342 35578 868 35588
rect 342 35512 352 35578
rect 858 35512 868 35578
rect 342 35502 868 35512
rect 970 35482 1500 35492
rect 970 35416 980 35482
rect 1490 35416 1500 35482
rect 970 35406 1500 35416
rect 342 35386 868 35396
rect 342 35320 352 35386
rect 858 35320 868 35386
rect 342 35310 868 35320
rect 970 35290 1500 35300
rect 970 35224 980 35290
rect 1490 35224 1500 35290
rect 970 35214 1500 35224
rect 342 35194 868 35204
rect 342 35128 352 35194
rect 858 35128 868 35194
rect 342 35118 868 35128
rect 970 35098 1500 35108
rect 970 35032 980 35098
rect 1490 35032 1500 35098
rect 970 35022 1500 35032
rect 342 35002 868 35012
rect 342 34936 352 35002
rect 858 34936 868 35002
rect 342 34926 868 34936
rect 970 34906 1500 34916
rect 970 34840 980 34906
rect 1490 34840 1500 34906
rect 970 34830 1500 34840
rect 342 34810 868 34820
rect 342 34744 352 34810
rect 858 34744 868 34810
rect 342 34734 868 34744
rect 970 34714 1500 34724
rect 970 34648 980 34714
rect 1490 34648 1500 34714
rect 970 34638 1500 34648
rect 342 34618 868 34628
rect 342 34552 352 34618
rect 858 34552 868 34618
rect 342 34542 868 34552
rect 970 34522 1500 34532
rect 970 34456 980 34522
rect 1490 34456 1500 34522
rect 970 34446 1500 34456
rect 342 34426 868 34436
rect 342 34360 352 34426
rect 858 34360 868 34426
rect 342 34350 868 34360
rect 970 34330 1500 34340
rect 970 34264 980 34330
rect 1490 34264 1500 34330
rect 970 34254 1500 34264
rect 342 34234 868 34244
rect 342 34168 352 34234
rect 858 34168 868 34234
rect 342 34158 868 34168
rect 970 34138 1500 34148
rect 970 34072 980 34138
rect 1490 34072 1500 34138
rect 970 34062 1500 34072
rect 342 34042 868 34052
rect 342 33976 352 34042
rect 858 33976 868 34042
rect 342 33966 868 33976
rect 970 33946 1500 33956
rect 970 33880 980 33946
rect 1490 33880 1500 33946
rect 970 33870 1500 33880
rect 342 33850 868 33860
rect 342 33784 352 33850
rect 858 33784 868 33850
rect 342 33774 868 33784
rect 970 33754 1500 33764
rect 970 33688 980 33754
rect 1490 33688 1500 33754
rect 970 33678 1500 33688
rect 342 33658 868 33668
rect 342 33592 352 33658
rect 858 33592 868 33658
rect 342 33582 868 33592
rect 970 33562 1500 33572
rect 970 33496 980 33562
rect 1490 33496 1500 33562
rect 970 33486 1500 33496
rect 342 33466 868 33476
rect 342 33400 352 33466
rect 858 33400 868 33466
rect 342 33390 868 33400
rect 970 33370 1500 33380
rect 970 33304 980 33370
rect 1490 33304 1500 33370
rect 970 33294 1500 33304
rect 342 33274 868 33284
rect 342 33208 352 33274
rect 858 33208 868 33274
rect 342 33198 868 33208
rect 970 33178 1500 33188
rect 970 33112 980 33178
rect 1490 33112 1500 33178
rect 970 33102 1500 33112
rect 342 33082 868 33092
rect 342 33016 352 33082
rect 858 33016 868 33082
rect 342 33006 868 33016
rect 970 32986 1500 32996
rect 970 32920 980 32986
rect 1490 32920 1500 32986
rect 970 32910 1500 32920
rect 342 32890 868 32900
rect 342 32824 352 32890
rect 858 32824 868 32890
rect 342 32814 868 32824
rect 970 32794 1500 32804
rect 970 32728 980 32794
rect 1490 32728 1500 32794
rect 970 32718 1500 32728
rect 342 32698 868 32708
rect 342 32632 352 32698
rect 858 32632 868 32698
rect 342 32622 868 32632
rect 970 32602 1500 32612
rect 970 32536 980 32602
rect 1490 32536 1500 32602
rect 970 32526 1500 32536
rect 342 32506 868 32516
rect 342 32440 352 32506
rect 858 32440 868 32506
rect 342 32430 868 32440
rect 970 32410 1500 32420
rect 970 32344 980 32410
rect 1490 32344 1500 32410
rect 970 32334 1500 32344
rect 342 32314 868 32324
rect 342 32248 352 32314
rect 858 32248 868 32314
rect 342 32238 868 32248
rect 970 32218 1500 32228
rect 970 32152 980 32218
rect 1490 32152 1500 32218
rect 970 32142 1500 32152
rect 342 32122 868 32132
rect 342 32056 352 32122
rect 858 32056 868 32122
rect 342 32046 868 32056
rect 970 32026 1500 32036
rect 970 31960 980 32026
rect 1490 31960 1500 32026
rect 970 31950 1500 31960
rect 342 31930 868 31940
rect 342 31864 352 31930
rect 858 31864 868 31930
rect 342 31854 868 31864
rect 970 31834 1500 31844
rect 970 31768 980 31834
rect 1490 31768 1500 31834
rect 970 31758 1500 31768
rect 342 31738 868 31748
rect 342 31672 352 31738
rect 858 31672 868 31738
rect 342 31662 868 31672
rect 970 31642 1500 31652
rect 970 31576 980 31642
rect 1490 31576 1500 31642
rect 970 31566 1500 31576
rect 342 31546 868 31556
rect 342 31480 352 31546
rect 858 31480 868 31546
rect 342 31470 868 31480
rect 970 31450 1500 31460
rect 970 31384 980 31450
rect 1490 31384 1500 31450
rect 970 31374 1500 31384
rect 342 31354 868 31364
rect 342 31288 352 31354
rect 858 31288 868 31354
rect 342 31278 868 31288
rect 970 31258 1500 31268
rect 970 31192 980 31258
rect 1490 31192 1500 31258
rect 970 31182 1500 31192
rect 342 31162 868 31172
rect 342 31096 352 31162
rect 858 31096 868 31162
rect 342 31086 868 31096
rect 970 31066 1500 31076
rect 970 31000 980 31066
rect 1490 31000 1500 31066
rect 970 30990 1500 31000
rect 342 30970 868 30980
rect 342 30904 352 30970
rect 858 30904 868 30970
rect 342 30894 868 30904
rect 970 30874 1500 30884
rect 970 30808 980 30874
rect 1490 30808 1500 30874
rect 970 30798 1500 30808
rect 342 30778 868 30788
rect 342 30712 352 30778
rect 858 30712 868 30778
rect 342 30702 868 30712
rect 970 30682 1500 30692
rect 970 30616 980 30682
rect 1490 30616 1500 30682
rect 970 30606 1500 30616
rect 342 30586 868 30596
rect 342 30520 352 30586
rect 858 30520 868 30586
rect 342 30510 868 30520
rect 970 30490 1500 30500
rect 970 30424 980 30490
rect 1490 30424 1500 30490
rect 970 30414 1500 30424
rect 342 30394 868 30404
rect 342 30328 352 30394
rect 858 30328 868 30394
rect 342 30318 868 30328
rect 970 30298 1500 30308
rect 970 30232 980 30298
rect 1490 30232 1500 30298
rect 970 30222 1500 30232
rect 342 30202 868 30212
rect 342 30136 352 30202
rect 858 30136 868 30202
rect 342 30126 868 30136
rect 970 30106 1500 30116
rect 970 30040 980 30106
rect 1490 30040 1500 30106
rect 970 30030 1500 30040
rect 342 30010 868 30020
rect 342 29944 352 30010
rect 858 29944 868 30010
rect 342 29934 868 29944
rect 970 29914 1500 29924
rect 970 29848 980 29914
rect 1490 29848 1500 29914
rect 970 29838 1500 29848
rect 342 29818 868 29828
rect 342 29752 352 29818
rect 858 29752 868 29818
rect 342 29742 868 29752
rect 970 29722 1500 29732
rect 970 29656 980 29722
rect 1490 29656 1500 29722
rect 970 29646 1500 29656
rect 342 29626 868 29636
rect 342 29560 352 29626
rect 858 29560 868 29626
rect 342 29550 868 29560
rect 970 29530 1500 29540
rect 970 29464 980 29530
rect 1490 29464 1500 29530
rect 970 29454 1500 29464
rect 342 29434 868 29444
rect 342 29368 352 29434
rect 858 29368 868 29434
rect 342 29358 868 29368
rect 970 29338 1500 29348
rect 970 29272 980 29338
rect 1490 29272 1500 29338
rect 970 29262 1500 29272
rect 342 29242 868 29252
rect 342 29176 352 29242
rect 858 29176 868 29242
rect 342 29166 868 29176
rect 970 29146 1500 29156
rect 970 29080 980 29146
rect 1490 29080 1500 29146
rect 970 29070 1500 29080
rect 342 29050 868 29060
rect 342 28984 352 29050
rect 858 28984 868 29050
rect 342 28974 868 28984
rect 970 28954 1500 28964
rect 970 28888 980 28954
rect 1490 28888 1500 28954
rect 970 28878 1500 28888
rect 342 28858 868 28868
rect 342 28792 352 28858
rect 858 28792 868 28858
rect 342 28782 868 28792
rect 970 28762 1500 28772
rect 970 28696 980 28762
rect 1490 28696 1500 28762
rect 970 28686 1500 28696
rect 342 28666 868 28676
rect 342 28600 352 28666
rect 858 28600 868 28666
rect 342 28590 868 28600
rect 970 28570 1500 28580
rect 970 28504 980 28570
rect 1490 28504 1500 28570
rect 970 28494 1500 28504
rect 342 28474 868 28484
rect 342 28408 352 28474
rect 858 28408 868 28474
rect 342 28398 868 28408
rect 970 28378 1500 28388
rect 970 28312 980 28378
rect 1490 28312 1500 28378
rect 970 28302 1500 28312
rect 342 28282 868 28292
rect 342 28216 352 28282
rect 858 28216 868 28282
rect 342 28206 868 28216
rect 970 28186 1500 28196
rect 970 28120 980 28186
rect 1490 28120 1500 28186
rect 970 28110 1500 28120
rect 342 28090 868 28100
rect 342 28024 352 28090
rect 858 28024 868 28090
rect 342 28014 868 28024
rect 970 27994 1500 28004
rect 970 27928 980 27994
rect 1490 27928 1500 27994
rect 970 27918 1500 27928
rect 342 27898 868 27908
rect 342 27832 352 27898
rect 858 27832 868 27898
rect 342 27822 868 27832
rect 970 27802 1500 27812
rect 970 27736 980 27802
rect 1490 27736 1500 27802
rect 970 27726 1500 27736
rect 342 27706 868 27716
rect 342 27640 352 27706
rect 858 27640 868 27706
rect 342 27630 868 27640
rect 970 27610 1500 27620
rect 970 27544 980 27610
rect 1490 27544 1500 27610
rect 970 27534 1500 27544
rect 342 27514 868 27524
rect 342 27448 352 27514
rect 858 27448 868 27514
rect 342 27438 868 27448
rect 970 27418 1500 27428
rect 970 27352 980 27418
rect 1490 27352 1500 27418
rect 970 27342 1500 27352
rect 342 27322 868 27332
rect 342 27256 352 27322
rect 858 27256 868 27322
rect 342 27246 868 27256
rect 970 27226 1500 27236
rect 970 27160 980 27226
rect 1490 27160 1500 27226
rect 970 27150 1500 27160
rect 342 27130 868 27140
rect 342 27064 352 27130
rect 858 27064 868 27130
rect 342 27054 868 27064
rect 970 27034 1500 27044
rect 970 26968 980 27034
rect 1490 26968 1500 27034
rect 970 26958 1500 26968
rect 342 26938 868 26948
rect 342 26872 352 26938
rect 858 26872 868 26938
rect 342 26862 868 26872
rect 970 26842 1500 26852
rect 970 26776 980 26842
rect 1490 26776 1500 26842
rect 970 26766 1500 26776
rect 342 26746 868 26756
rect 342 26680 352 26746
rect 858 26680 868 26746
rect 342 26670 868 26680
rect 970 26650 1500 26660
rect 970 26584 980 26650
rect 1490 26584 1500 26650
rect 970 26574 1500 26584
rect 342 26554 868 26564
rect 342 26488 352 26554
rect 858 26488 868 26554
rect 342 26478 868 26488
rect 970 26458 1500 26468
rect 970 26392 980 26458
rect 1490 26392 1500 26458
rect 970 26382 1500 26392
rect 342 26362 868 26372
rect 342 26296 352 26362
rect 858 26296 868 26362
rect 342 26286 868 26296
rect 970 26266 1500 26276
rect 970 26200 980 26266
rect 1490 26200 1500 26266
rect 970 26190 1500 26200
rect 342 26170 868 26180
rect 342 26104 352 26170
rect 858 26104 868 26170
rect 342 26094 868 26104
rect 970 26074 1500 26084
rect 970 26008 980 26074
rect 1490 26008 1500 26074
rect 970 25998 1500 26008
rect 342 25978 868 25988
rect 342 25912 352 25978
rect 858 25912 868 25978
rect 342 25902 868 25912
rect 970 25882 1500 25892
rect 970 25816 980 25882
rect 1490 25816 1500 25882
rect 970 25806 1500 25816
rect 342 25786 868 25796
rect 342 25720 352 25786
rect 858 25720 868 25786
rect 342 25710 868 25720
rect 970 25690 1500 25700
rect 970 25624 980 25690
rect 1490 25624 1500 25690
rect 970 25614 1500 25624
rect 342 25594 868 25604
rect 342 25528 352 25594
rect 858 25528 868 25594
rect 342 25518 868 25528
rect 970 25498 1500 25508
rect 970 25432 980 25498
rect 1490 25432 1500 25498
rect 970 25422 1500 25432
rect 342 25402 868 25412
rect 342 25336 352 25402
rect 858 25336 868 25402
rect 342 25326 868 25336
rect 970 25306 1500 25316
rect 970 25240 980 25306
rect 1490 25240 1500 25306
rect 970 25230 1500 25240
rect 342 25210 868 25220
rect 342 25144 352 25210
rect 858 25144 868 25210
rect 342 25134 868 25144
rect 970 25114 1500 25124
rect 970 25048 980 25114
rect 1490 25048 1500 25114
rect 970 25038 1500 25048
rect 342 25018 868 25028
rect 342 24952 352 25018
rect 858 24952 868 25018
rect 342 24942 868 24952
rect 970 24922 1500 24932
rect 970 24856 980 24922
rect 1490 24856 1500 24922
rect 970 24846 1500 24856
rect 342 24826 868 24836
rect 342 24760 352 24826
rect 858 24760 868 24826
rect 342 24750 868 24760
rect 970 24730 1500 24740
rect 970 24664 980 24730
rect 1490 24664 1500 24730
rect 970 24654 1500 24664
rect 342 24634 868 24644
rect 342 24568 352 24634
rect 858 24568 868 24634
rect 342 24558 868 24568
rect 970 24538 1500 24548
rect 970 24472 980 24538
rect 1490 24472 1500 24538
rect 970 24462 1500 24472
rect 342 24442 868 24452
rect 342 24376 352 24442
rect 858 24376 868 24442
rect 342 24366 868 24376
rect 970 24346 1500 24356
rect 970 24280 980 24346
rect 1490 24280 1500 24346
rect 970 24270 1500 24280
rect 342 24250 868 24260
rect 342 24184 352 24250
rect 858 24184 868 24250
rect 342 24174 868 24184
rect 970 24154 1500 24164
rect 970 24088 980 24154
rect 1490 24088 1500 24154
rect 970 24078 1500 24088
rect 342 24058 868 24068
rect 342 23992 352 24058
rect 858 23992 868 24058
rect 342 23982 868 23992
rect 970 23962 1500 23972
rect 970 23896 980 23962
rect 1490 23896 1500 23962
rect 970 23886 1500 23896
rect 342 23866 868 23876
rect 342 23800 352 23866
rect 858 23800 868 23866
rect 342 23790 868 23800
rect 970 23770 1500 23780
rect 970 23704 980 23770
rect 1490 23704 1500 23770
rect 970 23694 1500 23704
rect 342 23674 868 23684
rect 342 23608 352 23674
rect 858 23608 868 23674
rect 342 23598 868 23608
rect 970 23578 1500 23588
rect 970 23512 980 23578
rect 1490 23512 1500 23578
rect 970 23502 1500 23512
rect 342 23482 868 23492
rect 342 23416 352 23482
rect 858 23416 868 23482
rect 342 23406 868 23416
rect 970 23386 1500 23396
rect 970 23320 980 23386
rect 1490 23320 1500 23386
rect 970 23310 1500 23320
rect 342 23290 868 23300
rect 342 23224 352 23290
rect 858 23224 868 23290
rect 342 23214 868 23224
rect 970 23194 1500 23204
rect 970 23128 980 23194
rect 1490 23128 1500 23194
rect 970 23118 1500 23128
rect 342 23098 868 23108
rect 342 23032 352 23098
rect 858 23032 868 23098
rect 342 23022 868 23032
rect 340 22768 870 22778
rect 340 21976 870 21986
rect 342 21720 868 21730
rect 342 21654 352 21720
rect 858 21654 868 21720
rect 342 21644 868 21654
rect 970 21624 1500 21634
rect 970 21558 980 21624
rect 1490 21558 1500 21624
rect 970 21548 1500 21558
rect 342 21528 868 21538
rect 342 21462 352 21528
rect 858 21462 868 21528
rect 342 21452 868 21462
rect 970 21432 1500 21442
rect 970 21366 980 21432
rect 1490 21366 1500 21432
rect 970 21356 1500 21366
rect 342 21336 868 21346
rect 342 21270 352 21336
rect 858 21270 868 21336
rect 342 21260 868 21270
rect 970 21240 1500 21250
rect 970 21174 980 21240
rect 1490 21174 1500 21240
rect 970 21164 1500 21174
rect 342 21144 868 21154
rect 342 21078 352 21144
rect 858 21078 868 21144
rect 342 21068 868 21078
rect 970 21048 1500 21058
rect 970 20982 980 21048
rect 1490 20982 1500 21048
rect 970 20972 1500 20982
rect 342 20952 868 20962
rect 342 20886 352 20952
rect 858 20886 868 20952
rect 342 20876 868 20886
rect 970 20856 1500 20866
rect 970 20790 980 20856
rect 1490 20790 1500 20856
rect 970 20780 1500 20790
rect 342 20760 868 20770
rect 342 20694 352 20760
rect 858 20694 868 20760
rect 342 20684 868 20694
rect 970 20664 1500 20674
rect 970 20598 980 20664
rect 1490 20598 1500 20664
rect 970 20588 1500 20598
rect 342 20568 868 20578
rect 342 20502 352 20568
rect 858 20502 868 20568
rect 342 20492 868 20502
rect 970 20472 1500 20482
rect 970 20406 980 20472
rect 1490 20406 1500 20472
rect 970 20396 1500 20406
rect 342 20376 868 20386
rect 342 20310 352 20376
rect 858 20310 868 20376
rect 342 20300 868 20310
rect 970 20280 1500 20290
rect 970 20214 980 20280
rect 1490 20214 1500 20280
rect 970 20204 1500 20214
rect 342 20184 868 20194
rect 342 20118 352 20184
rect 858 20118 868 20184
rect 342 20108 868 20118
rect 970 20088 1500 20098
rect 970 20022 980 20088
rect 1490 20022 1500 20088
rect 970 20012 1500 20022
rect 342 19992 868 20002
rect 342 19926 352 19992
rect 858 19926 868 19992
rect 342 19916 868 19926
rect 970 19896 1500 19906
rect 970 19830 980 19896
rect 1490 19830 1500 19896
rect 970 19820 1500 19830
rect 342 19800 868 19810
rect 342 19734 352 19800
rect 858 19734 868 19800
rect 342 19724 868 19734
rect 970 19704 1500 19714
rect 970 19638 980 19704
rect 1490 19638 1500 19704
rect 970 19628 1500 19638
rect 342 19608 868 19618
rect 342 19542 352 19608
rect 858 19542 868 19608
rect 342 19532 868 19542
rect 970 19512 1500 19522
rect 970 19446 980 19512
rect 1490 19446 1500 19512
rect 970 19436 1500 19446
rect 342 19416 868 19426
rect 342 19350 352 19416
rect 858 19350 868 19416
rect 342 19340 868 19350
rect 970 19320 1500 19330
rect 970 19254 980 19320
rect 1490 19254 1500 19320
rect 970 19244 1500 19254
rect 342 19224 868 19234
rect 342 19158 352 19224
rect 858 19158 868 19224
rect 342 19148 868 19158
rect 970 19128 1500 19138
rect 970 19062 980 19128
rect 1490 19062 1500 19128
rect 970 19052 1500 19062
rect 342 19032 868 19042
rect 342 18966 352 19032
rect 858 18966 868 19032
rect 342 18956 868 18966
rect 970 18936 1500 18946
rect 970 18870 980 18936
rect 1490 18870 1500 18936
rect 970 18860 1500 18870
rect 342 18840 868 18850
rect 342 18774 352 18840
rect 858 18774 868 18840
rect 342 18764 868 18774
rect 970 18744 1500 18754
rect 970 18678 980 18744
rect 1490 18678 1500 18744
rect 970 18668 1500 18678
rect 342 18648 868 18658
rect 342 18582 352 18648
rect 858 18582 868 18648
rect 342 18572 868 18582
rect 970 18552 1500 18562
rect 970 18486 980 18552
rect 1490 18486 1500 18552
rect 970 18476 1500 18486
rect 342 18456 868 18466
rect 342 18390 352 18456
rect 858 18390 868 18456
rect 342 18380 868 18390
rect 970 18360 1500 18370
rect 970 18294 980 18360
rect 1490 18294 1500 18360
rect 970 18284 1500 18294
rect 342 18264 868 18274
rect 342 18198 352 18264
rect 858 18198 868 18264
rect 342 18188 868 18198
rect 970 18168 1500 18178
rect 970 18102 980 18168
rect 1490 18102 1500 18168
rect 970 18092 1500 18102
rect 342 18072 868 18082
rect 342 18006 352 18072
rect 858 18006 868 18072
rect 342 17996 868 18006
rect 970 17976 1500 17986
rect 970 17910 980 17976
rect 1490 17910 1500 17976
rect 970 17900 1500 17910
rect 342 17880 868 17890
rect 342 17814 352 17880
rect 858 17814 868 17880
rect 342 17804 868 17814
rect 970 17784 1500 17794
rect 970 17718 980 17784
rect 1490 17718 1500 17784
rect 970 17708 1500 17718
rect 342 17688 868 17698
rect 342 17622 352 17688
rect 858 17622 868 17688
rect 342 17612 868 17622
rect 970 17592 1500 17602
rect 970 17526 980 17592
rect 1490 17526 1500 17592
rect 970 17516 1500 17526
rect 342 17496 868 17506
rect 342 17430 352 17496
rect 858 17430 868 17496
rect 342 17420 868 17430
rect 970 17400 1500 17410
rect 970 17334 980 17400
rect 1490 17334 1500 17400
rect 970 17324 1500 17334
rect 342 17304 868 17314
rect 342 17238 352 17304
rect 858 17238 868 17304
rect 342 17228 868 17238
rect 970 17208 1500 17218
rect 970 17142 980 17208
rect 1490 17142 1500 17208
rect 970 17132 1500 17142
rect 342 17112 868 17122
rect 342 17046 352 17112
rect 858 17046 868 17112
rect 342 17036 868 17046
rect 970 17016 1500 17026
rect 970 16950 980 17016
rect 1490 16950 1500 17016
rect 970 16940 1500 16950
rect 342 16920 868 16930
rect 342 16854 352 16920
rect 858 16854 868 16920
rect 342 16844 868 16854
rect 970 16824 1500 16834
rect 970 16758 980 16824
rect 1490 16758 1500 16824
rect 970 16748 1500 16758
rect 342 16728 868 16738
rect 342 16662 352 16728
rect 858 16662 868 16728
rect 342 16652 868 16662
rect 970 16632 1500 16642
rect 970 16566 980 16632
rect 1490 16566 1500 16632
rect 970 16556 1500 16566
rect 342 16536 868 16546
rect 342 16470 352 16536
rect 858 16470 868 16536
rect 342 16460 868 16470
rect 970 16440 1500 16450
rect 970 16374 980 16440
rect 1490 16374 1500 16440
rect 970 16364 1500 16374
rect 342 16344 868 16354
rect 342 16278 352 16344
rect 858 16278 868 16344
rect 342 16268 868 16278
rect 970 16248 1500 16258
rect 970 16182 980 16248
rect 1490 16182 1500 16248
rect 970 16172 1500 16182
rect 342 16152 868 16162
rect 342 16086 352 16152
rect 858 16086 868 16152
rect 342 16076 868 16086
rect 970 16056 1500 16066
rect 970 15990 980 16056
rect 1490 15990 1500 16056
rect 970 15980 1500 15990
rect 342 15960 868 15970
rect 342 15894 352 15960
rect 858 15894 868 15960
rect 342 15884 868 15894
rect 970 15864 1500 15874
rect 970 15798 980 15864
rect 1490 15798 1500 15864
rect 970 15788 1500 15798
rect 342 15768 868 15778
rect 342 15702 352 15768
rect 858 15702 868 15768
rect 342 15692 868 15702
rect 970 15672 1500 15682
rect 970 15606 980 15672
rect 1490 15606 1500 15672
rect 970 15596 1500 15606
rect 342 15576 868 15586
rect 342 15510 352 15576
rect 858 15510 868 15576
rect 342 15500 868 15510
rect 970 15480 1500 15490
rect 970 15414 980 15480
rect 1490 15414 1500 15480
rect 970 15404 1500 15414
rect 342 15384 868 15394
rect 342 15318 352 15384
rect 858 15318 868 15384
rect 342 15308 868 15318
rect 970 15288 1500 15298
rect 970 15222 980 15288
rect 1490 15222 1500 15288
rect 970 15212 1500 15222
rect 342 15192 868 15202
rect 342 15126 352 15192
rect 858 15126 868 15192
rect 342 15116 868 15126
rect 970 15096 1500 15106
rect 970 15030 980 15096
rect 1490 15030 1500 15096
rect 970 15020 1500 15030
rect 342 15000 868 15010
rect 342 14934 352 15000
rect 858 14934 868 15000
rect 342 14924 868 14934
rect 970 14904 1500 14914
rect 970 14838 980 14904
rect 1490 14838 1500 14904
rect 970 14828 1500 14838
rect 342 14808 868 14818
rect 342 14742 352 14808
rect 858 14742 868 14808
rect 342 14732 868 14742
rect 970 14712 1500 14722
rect 970 14646 980 14712
rect 1490 14646 1500 14712
rect 970 14636 1500 14646
rect 342 14616 868 14626
rect 342 14550 352 14616
rect 858 14550 868 14616
rect 342 14540 868 14550
rect 970 14520 1500 14530
rect 970 14454 980 14520
rect 1490 14454 1500 14520
rect 970 14444 1500 14454
rect 342 14424 868 14434
rect 342 14358 352 14424
rect 858 14358 868 14424
rect 342 14348 868 14358
rect 970 14328 1500 14338
rect 970 14262 980 14328
rect 1490 14262 1500 14328
rect 970 14252 1500 14262
rect 342 14232 868 14242
rect 342 14166 352 14232
rect 858 14166 868 14232
rect 342 14156 868 14166
rect 970 14136 1500 14146
rect 970 14070 980 14136
rect 1490 14070 1500 14136
rect 970 14060 1500 14070
rect 342 14040 868 14050
rect 342 13974 352 14040
rect 858 13974 868 14040
rect 342 13964 868 13974
rect 970 13944 1500 13954
rect 970 13878 980 13944
rect 1490 13878 1500 13944
rect 970 13868 1500 13878
rect 342 13848 868 13858
rect 342 13782 352 13848
rect 858 13782 868 13848
rect 342 13772 868 13782
rect 970 13752 1500 13762
rect 970 13686 980 13752
rect 1490 13686 1500 13752
rect 970 13676 1500 13686
rect 342 13656 868 13666
rect 342 13590 352 13656
rect 858 13590 868 13656
rect 342 13580 868 13590
rect 970 13560 1500 13570
rect 970 13494 980 13560
rect 1490 13494 1500 13560
rect 970 13484 1500 13494
rect 342 13464 868 13474
rect 342 13398 352 13464
rect 858 13398 868 13464
rect 342 13388 868 13398
rect 970 13368 1500 13378
rect 970 13302 980 13368
rect 1490 13302 1500 13368
rect 970 13292 1500 13302
rect 342 13272 868 13282
rect 342 13206 352 13272
rect 858 13206 868 13272
rect 342 13196 868 13206
rect 970 13176 1500 13186
rect 970 13110 980 13176
rect 1490 13110 1500 13176
rect 970 13100 1500 13110
rect 342 13080 868 13090
rect 342 13014 352 13080
rect 858 13014 868 13080
rect 342 13004 868 13014
rect 970 12984 1500 12994
rect 970 12918 980 12984
rect 1490 12918 1500 12984
rect 970 12908 1500 12918
rect 342 12888 868 12898
rect 342 12822 352 12888
rect 858 12822 868 12888
rect 342 12812 868 12822
rect 970 12792 1500 12802
rect 970 12726 980 12792
rect 1490 12726 1500 12792
rect 970 12716 1500 12726
rect 342 12696 868 12706
rect 342 12630 352 12696
rect 858 12630 868 12696
rect 342 12620 868 12630
rect 970 12600 1500 12610
rect 970 12534 980 12600
rect 1490 12534 1500 12600
rect 970 12524 1500 12534
rect 342 12504 868 12514
rect 342 12438 352 12504
rect 858 12438 868 12504
rect 342 12428 868 12438
rect 970 12408 1500 12418
rect 970 12342 980 12408
rect 1490 12342 1500 12408
rect 970 12332 1500 12342
rect 342 12312 868 12322
rect 342 12246 352 12312
rect 858 12246 868 12312
rect 342 12236 868 12246
rect 970 12216 1500 12226
rect 970 12150 980 12216
rect 1490 12150 1500 12216
rect 970 12140 1500 12150
rect 342 12120 868 12130
rect 342 12054 352 12120
rect 858 12054 868 12120
rect 342 12044 868 12054
rect 970 12024 1500 12034
rect 970 11958 980 12024
rect 1490 11958 1500 12024
rect 970 11948 1500 11958
rect 342 11928 868 11938
rect 342 11862 352 11928
rect 858 11862 868 11928
rect 342 11852 868 11862
rect 970 11832 1500 11842
rect 970 11766 980 11832
rect 1490 11766 1500 11832
rect 970 11756 1500 11766
rect 342 11736 868 11746
rect 342 11670 352 11736
rect 858 11670 868 11736
rect 342 11660 868 11670
rect 970 11640 1500 11650
rect 970 11574 980 11640
rect 1490 11574 1500 11640
rect 970 11564 1500 11574
rect 342 11544 868 11554
rect 342 11478 352 11544
rect 858 11478 868 11544
rect 342 11468 868 11478
rect 970 11448 1500 11458
rect 970 11382 980 11448
rect 1490 11382 1500 11448
rect 970 11372 1500 11382
rect 342 11352 868 11362
rect 342 11286 352 11352
rect 858 11286 868 11352
rect 342 11276 868 11286
rect 970 11256 1500 11266
rect 970 11190 980 11256
rect 1490 11190 1500 11256
rect 970 11180 1500 11190
rect 342 11160 868 11170
rect 342 11094 352 11160
rect 858 11094 868 11160
rect 342 11084 868 11094
rect 970 11064 1500 11074
rect 970 10998 980 11064
rect 1490 10998 1500 11064
rect 970 10988 1500 10998
rect 342 10968 868 10978
rect 342 10902 352 10968
rect 858 10902 868 10968
rect 342 10892 868 10902
rect 970 10872 1500 10882
rect 970 10806 980 10872
rect 1490 10806 1500 10872
rect 970 10796 1500 10806
rect 342 10776 868 10786
rect 342 10710 352 10776
rect 858 10710 868 10776
rect 342 10700 868 10710
rect 970 10680 1500 10690
rect 970 10614 980 10680
rect 1490 10614 1500 10680
rect 970 10604 1500 10614
rect 342 10584 868 10594
rect 342 10518 352 10584
rect 858 10518 868 10584
rect 342 10508 868 10518
rect 970 10488 1500 10498
rect 970 10422 980 10488
rect 1490 10422 1500 10488
rect 970 10412 1500 10422
rect 342 10392 868 10402
rect 342 10326 352 10392
rect 858 10326 868 10392
rect 342 10316 868 10326
rect 970 10296 1500 10306
rect 970 10230 980 10296
rect 1490 10230 1500 10296
rect 970 10220 1500 10230
rect 342 10200 868 10210
rect 342 10134 352 10200
rect 858 10134 868 10200
rect 342 10124 868 10134
rect 970 10104 1500 10114
rect 970 10038 980 10104
rect 1490 10038 1500 10104
rect 970 10028 1500 10038
rect 342 10008 868 10018
rect 342 9942 352 10008
rect 858 9942 868 10008
rect 342 9932 868 9942
rect 970 9912 1500 9922
rect 970 9846 980 9912
rect 1490 9846 1500 9912
rect 970 9836 1500 9846
rect 342 9816 868 9826
rect 342 9750 352 9816
rect 858 9750 868 9816
rect 342 9740 868 9750
rect 970 9720 1500 9730
rect 970 9654 980 9720
rect 1490 9654 1500 9720
rect 970 9644 1500 9654
rect 342 9624 868 9634
rect 342 9558 352 9624
rect 858 9558 868 9624
rect 342 9548 868 9558
rect 970 9528 1500 9538
rect 970 9462 980 9528
rect 1490 9462 1500 9528
rect 970 9452 1500 9462
rect 342 9432 868 9442
rect 342 9366 352 9432
rect 858 9366 868 9432
rect 342 9356 868 9366
rect 970 9336 1500 9346
rect 970 9270 980 9336
rect 1490 9270 1500 9336
rect 970 9260 1500 9270
rect 342 9240 868 9250
rect 342 9174 352 9240
rect 858 9174 868 9240
rect 342 9164 868 9174
rect 970 9144 1500 9154
rect 970 9078 980 9144
rect 1490 9078 1500 9144
rect 970 9068 1500 9078
rect 342 9048 868 9058
rect 342 8982 352 9048
rect 858 8982 868 9048
rect 342 8972 868 8982
rect 970 8952 1500 8962
rect 970 8886 980 8952
rect 1490 8886 1500 8952
rect 970 8876 1500 8886
rect 342 8856 868 8866
rect 342 8790 352 8856
rect 858 8790 868 8856
rect 342 8780 868 8790
rect 970 8760 1500 8770
rect 970 8694 980 8760
rect 1490 8694 1500 8760
rect 970 8684 1500 8694
rect 342 8664 868 8674
rect 342 8598 352 8664
rect 858 8598 868 8664
rect 342 8588 868 8598
rect 970 8568 1500 8578
rect 970 8502 980 8568
rect 1490 8502 1500 8568
rect 970 8492 1500 8502
rect 342 8472 868 8482
rect 342 8406 352 8472
rect 858 8406 868 8472
rect 342 8396 868 8406
rect 970 8376 1500 8386
rect 970 8310 980 8376
rect 1490 8310 1500 8376
rect 970 8300 1500 8310
rect 342 8280 868 8290
rect 342 8214 352 8280
rect 858 8214 868 8280
rect 342 8204 868 8214
rect 970 8184 1500 8194
rect 970 8118 980 8184
rect 1490 8118 1500 8184
rect 970 8108 1500 8118
rect 342 8088 868 8098
rect 342 8022 352 8088
rect 858 8022 868 8088
rect 342 8012 868 8022
rect 970 7992 1500 8002
rect 970 7926 980 7992
rect 1490 7926 1500 7992
rect 970 7916 1500 7926
rect 342 7896 868 7906
rect 342 7830 352 7896
rect 858 7830 868 7896
rect 342 7820 868 7830
rect 970 7800 1500 7810
rect 970 7734 980 7800
rect 1490 7734 1500 7800
rect 970 7724 1500 7734
rect 342 7704 868 7714
rect 342 7638 352 7704
rect 858 7638 868 7704
rect 342 7628 868 7638
rect 970 7608 1500 7618
rect 970 7542 980 7608
rect 1490 7542 1500 7608
rect 970 7532 1500 7542
rect 342 7512 868 7522
rect 342 7446 352 7512
rect 858 7446 868 7512
rect 342 7436 868 7446
rect 970 7416 1500 7426
rect 970 7350 980 7416
rect 1490 7350 1500 7416
rect 970 7340 1500 7350
rect 342 7320 868 7330
rect 342 7254 352 7320
rect 858 7254 868 7320
rect 342 7244 868 7254
rect 970 7224 1500 7234
rect 970 7158 980 7224
rect 1490 7158 1500 7224
rect 970 7148 1500 7158
rect 342 7128 868 7138
rect 342 7062 352 7128
rect 858 7062 868 7128
rect 342 7052 868 7062
rect 970 7032 1500 7042
rect 970 6966 980 7032
rect 1490 6966 1500 7032
rect 970 6956 1500 6966
rect 342 6936 868 6946
rect 342 6870 352 6936
rect 858 6870 868 6936
rect 342 6860 868 6870
rect 970 6840 1500 6850
rect 970 6774 980 6840
rect 1490 6774 1500 6840
rect 970 6764 1500 6774
rect 342 6744 868 6754
rect 342 6678 352 6744
rect 858 6678 868 6744
rect 342 6668 868 6678
rect 970 6648 1500 6658
rect 970 6582 980 6648
rect 1490 6582 1500 6648
rect 970 6572 1500 6582
rect 342 6552 868 6562
rect 342 6486 352 6552
rect 858 6486 868 6552
rect 342 6476 868 6486
rect 970 6456 1500 6466
rect 970 6390 980 6456
rect 1490 6390 1500 6456
rect 970 6380 1500 6390
rect 342 6360 868 6370
rect 342 6294 352 6360
rect 858 6294 868 6360
rect 342 6284 868 6294
rect 970 6264 1500 6274
rect 970 6198 980 6264
rect 1490 6198 1500 6264
rect 970 6188 1500 6198
rect 342 6168 868 6178
rect 342 6102 352 6168
rect 858 6102 868 6168
rect 342 6092 868 6102
rect 970 6072 1500 6082
rect 970 6006 980 6072
rect 1490 6006 1500 6072
rect 970 5996 1500 6006
rect 342 5976 868 5986
rect 342 5910 352 5976
rect 858 5910 868 5976
rect 342 5900 868 5910
rect 970 5880 1500 5890
rect 970 5814 980 5880
rect 1490 5814 1500 5880
rect 970 5804 1500 5814
rect 342 5784 868 5794
rect 342 5718 352 5784
rect 858 5718 868 5784
rect 342 5708 868 5718
rect 970 5688 1500 5698
rect 970 5622 980 5688
rect 1490 5622 1500 5688
rect 970 5612 1500 5622
rect 342 5592 868 5602
rect 342 5526 352 5592
rect 858 5526 868 5592
rect 342 5516 868 5526
rect 970 5496 1500 5506
rect 970 5430 980 5496
rect 1490 5430 1500 5496
rect 970 5420 1500 5430
rect 342 5400 868 5410
rect 342 5334 352 5400
rect 858 5334 868 5400
rect 342 5324 868 5334
rect 970 5304 1500 5314
rect 970 5238 980 5304
rect 1490 5238 1500 5304
rect 970 5228 1500 5238
rect 342 5208 868 5218
rect 342 5142 352 5208
rect 858 5142 868 5208
rect 342 5132 868 5142
rect 970 5112 1500 5122
rect 970 5046 980 5112
rect 1490 5046 1500 5112
rect 970 5036 1500 5046
rect 342 5016 868 5026
rect 342 4950 352 5016
rect 858 4950 868 5016
rect 342 4940 868 4950
rect 970 4920 1500 4930
rect 970 4854 980 4920
rect 1490 4854 1500 4920
rect 970 4844 1500 4854
rect 342 4824 868 4834
rect 342 4758 352 4824
rect 858 4758 868 4824
rect 342 4748 868 4758
rect 970 4728 1500 4738
rect 970 4662 980 4728
rect 1490 4662 1500 4728
rect 970 4652 1500 4662
rect 342 4632 868 4642
rect 342 4566 352 4632
rect 858 4566 868 4632
rect 342 4556 868 4566
rect 970 4536 1500 4546
rect 970 4470 980 4536
rect 1490 4470 1500 4536
rect 970 4460 1500 4470
rect 342 4440 868 4450
rect 342 4374 352 4440
rect 858 4374 868 4440
rect 342 4364 868 4374
rect 970 4344 1500 4354
rect 970 4278 980 4344
rect 1490 4278 1500 4344
rect 970 4268 1500 4278
rect 342 4248 868 4258
rect 342 4182 352 4248
rect 858 4182 868 4248
rect 342 4172 868 4182
rect 970 4152 1500 4162
rect 970 4086 980 4152
rect 1490 4086 1500 4152
rect 970 4076 1500 4086
rect 342 4056 868 4066
rect 342 3990 352 4056
rect 858 3990 868 4056
rect 342 3980 868 3990
rect 970 3960 1500 3970
rect 970 3894 980 3960
rect 1490 3894 1500 3960
rect 970 3884 1500 3894
rect 342 3864 868 3874
rect 342 3798 352 3864
rect 858 3798 868 3864
rect 342 3788 868 3798
rect 970 3768 1500 3778
rect 970 3702 980 3768
rect 1490 3702 1500 3768
rect 970 3692 1500 3702
rect 342 3672 868 3682
rect 342 3606 352 3672
rect 858 3606 868 3672
rect 342 3596 868 3606
rect 970 3576 1500 3586
rect 970 3510 980 3576
rect 1490 3510 1500 3576
rect 970 3500 1500 3510
rect 342 3480 868 3490
rect 342 3414 352 3480
rect 858 3414 868 3480
rect 342 3404 868 3414
rect 970 3384 1500 3394
rect 970 3318 980 3384
rect 1490 3318 1500 3384
rect 970 3308 1500 3318
rect 342 3288 868 3298
rect 342 3222 352 3288
rect 858 3222 868 3288
rect 342 3212 868 3222
rect 970 3192 1500 3202
rect 970 3126 980 3192
rect 1490 3126 1500 3192
rect 970 3116 1500 3126
rect 342 3096 868 3106
rect 342 3030 352 3096
rect 858 3030 868 3096
rect 342 3020 868 3030
rect 970 3000 1500 3010
rect 970 2934 980 3000
rect 1490 2934 1500 3000
rect 970 2924 1500 2934
rect 342 2904 868 2914
rect 342 2838 352 2904
rect 858 2838 868 2904
rect 342 2828 868 2838
rect 970 2808 1500 2818
rect 970 2742 980 2808
rect 1490 2742 1500 2808
rect 970 2732 1500 2742
rect 342 2712 868 2722
rect 342 2646 352 2712
rect 858 2646 868 2712
rect 342 2636 868 2646
rect 970 2616 1500 2626
rect 970 2550 980 2616
rect 1490 2550 1500 2616
rect 970 2540 1500 2550
rect 342 2520 868 2530
rect 342 2454 352 2520
rect 858 2454 868 2520
rect 342 2444 868 2454
rect 970 2424 1500 2434
rect 970 2358 980 2424
rect 1490 2358 1500 2424
rect 970 2348 1500 2358
rect 342 2328 868 2338
rect 342 2262 352 2328
rect 858 2262 868 2328
rect 342 2252 868 2262
rect 970 2232 1500 2242
rect 970 2166 980 2232
rect 1490 2166 1500 2232
rect 970 2156 1500 2166
rect 342 2136 868 2146
rect 342 2070 352 2136
rect 858 2070 868 2136
rect 342 2060 868 2070
rect 970 2040 1500 2050
rect 970 1974 980 2040
rect 1490 1974 1500 2040
rect 970 1964 1500 1974
rect 342 1944 868 1954
rect 342 1878 352 1944
rect 858 1878 868 1944
rect 342 1868 868 1878
rect 970 1848 1500 1858
rect 970 1782 980 1848
rect 1490 1782 1500 1848
rect 970 1772 1500 1782
rect 342 1752 868 1762
rect 342 1686 352 1752
rect 858 1686 868 1752
rect 342 1676 868 1686
rect 970 1656 1500 1666
rect 970 1590 980 1656
rect 1490 1590 1500 1656
rect 970 1580 1500 1590
rect 342 1560 868 1570
rect 342 1494 352 1560
rect 858 1494 868 1560
rect 342 1484 868 1494
rect 970 1464 1500 1474
rect 970 1398 980 1464
rect 1490 1398 1500 1464
rect 970 1388 1500 1398
rect 342 1368 868 1378
rect 342 1302 352 1368
rect 858 1302 868 1368
rect 342 1292 868 1302
rect 970 1272 1500 1282
rect 970 1206 980 1272
rect 1490 1206 1500 1272
rect 970 1196 1500 1206
rect 342 1176 868 1186
rect 342 1110 352 1176
rect 858 1110 868 1176
rect 342 1100 868 1110
rect 970 1080 1500 1090
rect 970 1014 980 1080
rect 1490 1014 1500 1080
rect 970 1004 1500 1014
rect 342 984 868 994
rect 342 918 352 984
rect 858 918 868 984
rect 342 908 868 918
rect 970 888 1500 898
rect 970 822 980 888
rect 1490 822 1500 888
rect 970 812 1500 822
rect 342 792 868 802
rect 342 726 352 792
rect 858 726 868 792
rect 342 716 868 726
rect 970 696 1500 706
rect 970 630 980 696
rect 1490 630 1500 696
rect 970 620 1500 630
rect 342 600 868 610
rect 342 534 352 600
rect 858 534 868 600
rect 342 524 868 534
<< via2 >>
rect 132 45126 1706 45136
rect 132 45072 1706 45126
rect 132 45062 1706 45072
rect 352 44152 858 44218
rect 980 44056 1490 44122
rect 352 43960 858 44026
rect 980 43864 1490 43930
rect 352 43768 858 43834
rect 980 43672 1490 43738
rect 352 43576 858 43642
rect 980 43480 1490 43546
rect 352 43384 858 43450
rect 980 43288 1490 43354
rect 352 43192 858 43258
rect 980 43096 1490 43162
rect 352 43000 858 43066
rect 980 42904 1490 42970
rect 352 42808 858 42874
rect 980 42712 1490 42778
rect 352 42616 858 42682
rect 980 42520 1490 42586
rect 352 42424 858 42490
rect 980 42328 1490 42394
rect 352 42232 858 42298
rect 980 42136 1490 42202
rect 352 42040 858 42106
rect 980 41944 1490 42010
rect 352 41848 858 41914
rect 980 41752 1490 41818
rect 352 41656 858 41722
rect 980 41560 1490 41626
rect 352 41464 858 41530
rect 980 41368 1490 41434
rect 352 41272 858 41338
rect 980 41176 1490 41242
rect 352 41080 858 41146
rect 980 40984 1490 41050
rect 352 40888 858 40954
rect 980 40792 1490 40858
rect 352 40696 858 40762
rect 980 40600 1490 40666
rect 352 40504 858 40570
rect 980 40408 1490 40474
rect 352 40312 858 40378
rect 980 40216 1490 40282
rect 352 40120 858 40186
rect 980 40024 1490 40090
rect 352 39928 858 39994
rect 980 39832 1490 39898
rect 352 39736 858 39802
rect 980 39640 1490 39706
rect 352 39544 858 39610
rect 980 39448 1490 39514
rect 352 39352 858 39418
rect 980 39256 1490 39322
rect 352 39160 858 39226
rect 980 39064 1490 39130
rect 352 38968 858 39034
rect 980 38872 1490 38938
rect 352 38776 858 38842
rect 980 38680 1490 38746
rect 352 38584 858 38650
rect 980 38488 1490 38554
rect 352 38392 858 38458
rect 980 38296 1490 38362
rect 352 38200 858 38266
rect 980 38104 1490 38170
rect 352 38008 858 38074
rect 980 37912 1490 37978
rect 352 37816 858 37882
rect 980 37720 1490 37786
rect 352 37624 858 37690
rect 980 37528 1490 37594
rect 352 37432 858 37498
rect 980 37336 1490 37402
rect 352 37240 858 37306
rect 980 37144 1490 37210
rect 352 37048 858 37114
rect 980 36952 1490 37018
rect 352 36856 858 36922
rect 980 36760 1490 36826
rect 352 36664 858 36730
rect 980 36568 1490 36634
rect 352 36472 858 36538
rect 980 36376 1490 36442
rect 352 36280 858 36346
rect 980 36184 1490 36250
rect 352 36088 858 36154
rect 980 35992 1490 36058
rect 352 35896 858 35962
rect 980 35800 1490 35866
rect 352 35704 858 35770
rect 980 35608 1490 35674
rect 352 35512 858 35578
rect 980 35416 1490 35482
rect 352 35320 858 35386
rect 980 35224 1490 35290
rect 352 35128 858 35194
rect 980 35032 1490 35098
rect 352 34936 858 35002
rect 980 34840 1490 34906
rect 352 34744 858 34810
rect 980 34648 1490 34714
rect 352 34552 858 34618
rect 980 34456 1490 34522
rect 352 34360 858 34426
rect 980 34264 1490 34330
rect 352 34168 858 34234
rect 980 34072 1490 34138
rect 352 33976 858 34042
rect 980 33880 1490 33946
rect 352 33784 858 33850
rect 980 33688 1490 33754
rect 352 33592 858 33658
rect 980 33496 1490 33562
rect 352 33400 858 33466
rect 980 33304 1490 33370
rect 352 33208 858 33274
rect 980 33112 1490 33178
rect 352 33016 858 33082
rect 980 32920 1490 32986
rect 352 32824 858 32890
rect 980 32728 1490 32794
rect 352 32632 858 32698
rect 980 32536 1490 32602
rect 352 32440 858 32506
rect 980 32344 1490 32410
rect 352 32248 858 32314
rect 980 32152 1490 32218
rect 352 32056 858 32122
rect 980 31960 1490 32026
rect 352 31864 858 31930
rect 980 31768 1490 31834
rect 352 31672 858 31738
rect 980 31576 1490 31642
rect 352 31480 858 31546
rect 980 31384 1490 31450
rect 352 31288 858 31354
rect 980 31192 1490 31258
rect 352 31096 858 31162
rect 980 31000 1490 31066
rect 352 30904 858 30970
rect 980 30808 1490 30874
rect 352 30712 858 30778
rect 980 30616 1490 30682
rect 352 30520 858 30586
rect 980 30424 1490 30490
rect 352 30328 858 30394
rect 980 30232 1490 30298
rect 352 30136 858 30202
rect 980 30040 1490 30106
rect 352 29944 858 30010
rect 980 29848 1490 29914
rect 352 29752 858 29818
rect 980 29656 1490 29722
rect 352 29560 858 29626
rect 980 29464 1490 29530
rect 352 29368 858 29434
rect 980 29272 1490 29338
rect 352 29176 858 29242
rect 980 29080 1490 29146
rect 352 28984 858 29050
rect 980 28888 1490 28954
rect 352 28792 858 28858
rect 980 28696 1490 28762
rect 352 28600 858 28666
rect 980 28504 1490 28570
rect 352 28408 858 28474
rect 980 28312 1490 28378
rect 352 28216 858 28282
rect 980 28120 1490 28186
rect 352 28024 858 28090
rect 980 27928 1490 27994
rect 352 27832 858 27898
rect 980 27736 1490 27802
rect 352 27640 858 27706
rect 980 27544 1490 27610
rect 352 27448 858 27514
rect 980 27352 1490 27418
rect 352 27256 858 27322
rect 980 27160 1490 27226
rect 352 27064 858 27130
rect 980 26968 1490 27034
rect 352 26872 858 26938
rect 980 26776 1490 26842
rect 352 26680 858 26746
rect 980 26584 1490 26650
rect 352 26488 858 26554
rect 980 26392 1490 26458
rect 352 26296 858 26362
rect 980 26200 1490 26266
rect 352 26104 858 26170
rect 980 26008 1490 26074
rect 352 25912 858 25978
rect 980 25816 1490 25882
rect 352 25720 858 25786
rect 980 25624 1490 25690
rect 352 25528 858 25594
rect 980 25432 1490 25498
rect 352 25336 858 25402
rect 980 25240 1490 25306
rect 352 25144 858 25210
rect 980 25048 1490 25114
rect 352 24952 858 25018
rect 980 24856 1490 24922
rect 352 24760 858 24826
rect 980 24664 1490 24730
rect 352 24568 858 24634
rect 980 24472 1490 24538
rect 352 24376 858 24442
rect 980 24280 1490 24346
rect 352 24184 858 24250
rect 980 24088 1490 24154
rect 352 23992 858 24058
rect 980 23896 1490 23962
rect 352 23800 858 23866
rect 980 23704 1490 23770
rect 352 23608 858 23674
rect 980 23512 1490 23578
rect 352 23416 858 23482
rect 980 23320 1490 23386
rect 352 23224 858 23290
rect 980 23128 1490 23194
rect 352 23032 858 23098
rect 340 21986 870 22768
rect 352 21654 858 21720
rect 980 21558 1490 21624
rect 352 21462 858 21528
rect 980 21366 1490 21432
rect 352 21270 858 21336
rect 980 21174 1490 21240
rect 352 21078 858 21144
rect 980 20982 1490 21048
rect 352 20886 858 20952
rect 980 20790 1490 20856
rect 352 20694 858 20760
rect 980 20598 1490 20664
rect 352 20502 858 20568
rect 980 20406 1490 20472
rect 352 20310 858 20376
rect 980 20214 1490 20280
rect 352 20118 858 20184
rect 980 20022 1490 20088
rect 352 19926 858 19992
rect 980 19830 1490 19896
rect 352 19734 858 19800
rect 980 19638 1490 19704
rect 352 19542 858 19608
rect 980 19446 1490 19512
rect 352 19350 858 19416
rect 980 19254 1490 19320
rect 352 19158 858 19224
rect 980 19062 1490 19128
rect 352 18966 858 19032
rect 980 18870 1490 18936
rect 352 18774 858 18840
rect 980 18678 1490 18744
rect 352 18582 858 18648
rect 980 18486 1490 18552
rect 352 18390 858 18456
rect 980 18294 1490 18360
rect 352 18198 858 18264
rect 980 18102 1490 18168
rect 352 18006 858 18072
rect 980 17910 1490 17976
rect 352 17814 858 17880
rect 980 17718 1490 17784
rect 352 17622 858 17688
rect 980 17526 1490 17592
rect 352 17430 858 17496
rect 980 17334 1490 17400
rect 352 17238 858 17304
rect 980 17142 1490 17208
rect 352 17046 858 17112
rect 980 16950 1490 17016
rect 352 16854 858 16920
rect 980 16758 1490 16824
rect 352 16662 858 16728
rect 980 16566 1490 16632
rect 352 16470 858 16536
rect 980 16374 1490 16440
rect 352 16278 858 16344
rect 980 16182 1490 16248
rect 352 16086 858 16152
rect 980 15990 1490 16056
rect 352 15894 858 15960
rect 980 15798 1490 15864
rect 352 15702 858 15768
rect 980 15606 1490 15672
rect 352 15510 858 15576
rect 980 15414 1490 15480
rect 352 15318 858 15384
rect 980 15222 1490 15288
rect 352 15126 858 15192
rect 980 15030 1490 15096
rect 352 14934 858 15000
rect 980 14838 1490 14904
rect 352 14742 858 14808
rect 980 14646 1490 14712
rect 352 14550 858 14616
rect 980 14454 1490 14520
rect 352 14358 858 14424
rect 980 14262 1490 14328
rect 352 14166 858 14232
rect 980 14070 1490 14136
rect 352 13974 858 14040
rect 980 13878 1490 13944
rect 352 13782 858 13848
rect 980 13686 1490 13752
rect 352 13590 858 13656
rect 980 13494 1490 13560
rect 352 13398 858 13464
rect 980 13302 1490 13368
rect 352 13206 858 13272
rect 980 13110 1490 13176
rect 352 13014 858 13080
rect 980 12918 1490 12984
rect 352 12822 858 12888
rect 980 12726 1490 12792
rect 352 12630 858 12696
rect 980 12534 1490 12600
rect 352 12438 858 12504
rect 980 12342 1490 12408
rect 352 12246 858 12312
rect 980 12150 1490 12216
rect 352 12054 858 12120
rect 980 11958 1490 12024
rect 352 11862 858 11928
rect 980 11766 1490 11832
rect 352 11670 858 11736
rect 980 11574 1490 11640
rect 352 11478 858 11544
rect 980 11382 1490 11448
rect 352 11286 858 11352
rect 980 11190 1490 11256
rect 352 11094 858 11160
rect 980 10998 1490 11064
rect 352 10902 858 10968
rect 980 10806 1490 10872
rect 352 10710 858 10776
rect 980 10614 1490 10680
rect 352 10518 858 10584
rect 980 10422 1490 10488
rect 352 10326 858 10392
rect 980 10230 1490 10296
rect 352 10134 858 10200
rect 980 10038 1490 10104
rect 352 9942 858 10008
rect 980 9846 1490 9912
rect 352 9750 858 9816
rect 980 9654 1490 9720
rect 352 9558 858 9624
rect 980 9462 1490 9528
rect 352 9366 858 9432
rect 980 9270 1490 9336
rect 352 9174 858 9240
rect 980 9078 1490 9144
rect 352 8982 858 9048
rect 980 8886 1490 8952
rect 352 8790 858 8856
rect 980 8694 1490 8760
rect 352 8598 858 8664
rect 980 8502 1490 8568
rect 352 8406 858 8472
rect 980 8310 1490 8376
rect 352 8214 858 8280
rect 980 8118 1490 8184
rect 352 8022 858 8088
rect 980 7926 1490 7992
rect 352 7830 858 7896
rect 980 7734 1490 7800
rect 352 7638 858 7704
rect 980 7542 1490 7608
rect 352 7446 858 7512
rect 980 7350 1490 7416
rect 352 7254 858 7320
rect 980 7158 1490 7224
rect 352 7062 858 7128
rect 980 6966 1490 7032
rect 352 6870 858 6936
rect 980 6774 1490 6840
rect 352 6678 858 6744
rect 980 6582 1490 6648
rect 352 6486 858 6552
rect 980 6390 1490 6456
rect 352 6294 858 6360
rect 980 6198 1490 6264
rect 352 6102 858 6168
rect 980 6006 1490 6072
rect 352 5910 858 5976
rect 980 5814 1490 5880
rect 352 5718 858 5784
rect 980 5622 1490 5688
rect 352 5526 858 5592
rect 980 5430 1490 5496
rect 352 5334 858 5400
rect 980 5238 1490 5304
rect 352 5142 858 5208
rect 980 5046 1490 5112
rect 352 4950 858 5016
rect 980 4854 1490 4920
rect 352 4758 858 4824
rect 980 4662 1490 4728
rect 352 4566 858 4632
rect 980 4470 1490 4536
rect 352 4374 858 4440
rect 980 4278 1490 4344
rect 352 4182 858 4248
rect 980 4086 1490 4152
rect 352 3990 858 4056
rect 980 3894 1490 3960
rect 352 3798 858 3864
rect 980 3702 1490 3768
rect 352 3606 858 3672
rect 980 3510 1490 3576
rect 352 3414 858 3480
rect 980 3318 1490 3384
rect 352 3222 858 3288
rect 980 3126 1490 3192
rect 352 3030 858 3096
rect 980 2934 1490 3000
rect 352 2838 858 2904
rect 980 2742 1490 2808
rect 352 2646 858 2712
rect 980 2550 1490 2616
rect 352 2454 858 2520
rect 980 2358 1490 2424
rect 352 2262 858 2328
rect 980 2166 1490 2232
rect 352 2070 858 2136
rect 980 1974 1490 2040
rect 352 1878 858 1944
rect 980 1782 1490 1848
rect 352 1686 858 1752
rect 980 1590 1490 1656
rect 352 1494 858 1560
rect 980 1398 1490 1464
rect 352 1302 858 1368
rect 980 1206 1490 1272
rect 352 1110 858 1176
rect 980 1014 1490 1080
rect 352 918 858 984
rect 980 822 1490 888
rect 352 726 858 792
rect 980 630 1490 696
rect 352 534 858 600
<< metal3 >>
rect 122 45136 1716 45141
rect 122 45062 132 45136
rect 1706 45062 1716 45136
rect 122 45057 1716 45062
rect 342 44218 868 44228
rect 342 44152 352 44218
rect 858 44152 868 44218
rect 342 44142 868 44152
rect 970 44122 1500 44132
rect 970 44056 980 44122
rect 1490 44056 1500 44122
rect 970 44046 1500 44056
rect 342 44026 868 44036
rect 342 43960 352 44026
rect 858 43960 868 44026
rect 342 43950 868 43960
rect 970 43930 1500 43940
rect 970 43864 980 43930
rect 1490 43864 1500 43930
rect 970 43854 1500 43864
rect 342 43834 868 43844
rect 342 43768 352 43834
rect 858 43768 868 43834
rect 342 43758 868 43768
rect 970 43738 1500 43748
rect 970 43672 980 43738
rect 1490 43672 1500 43738
rect 970 43662 1500 43672
rect 342 43642 868 43652
rect 342 43576 352 43642
rect 858 43576 868 43642
rect 342 43566 868 43576
rect 970 43546 1500 43556
rect 970 43480 980 43546
rect 1490 43480 1500 43546
rect 970 43470 1500 43480
rect 342 43450 868 43460
rect 342 43384 352 43450
rect 858 43384 868 43450
rect 342 43374 868 43384
rect 970 43354 1500 43364
rect 970 43288 980 43354
rect 1490 43288 1500 43354
rect 970 43278 1500 43288
rect 342 43258 868 43268
rect 342 43192 352 43258
rect 858 43192 868 43258
rect 342 43182 868 43192
rect 970 43162 1500 43172
rect 970 43096 980 43162
rect 1490 43096 1500 43162
rect 970 43086 1500 43096
rect 342 43066 868 43076
rect 342 43000 352 43066
rect 858 43000 868 43066
rect 342 42990 868 43000
rect 970 42970 1500 42980
rect 970 42904 980 42970
rect 1490 42904 1500 42970
rect 970 42894 1500 42904
rect 342 42874 868 42884
rect 342 42808 352 42874
rect 858 42808 868 42874
rect 342 42798 868 42808
rect 970 42778 1500 42788
rect 970 42712 980 42778
rect 1490 42712 1500 42778
rect 970 42702 1500 42712
rect 342 42682 868 42692
rect 342 42616 352 42682
rect 858 42616 868 42682
rect 342 42606 868 42616
rect 970 42586 1500 42596
rect 970 42520 980 42586
rect 1490 42520 1500 42586
rect 970 42510 1500 42520
rect 342 42490 868 42500
rect 342 42424 352 42490
rect 858 42424 868 42490
rect 342 42414 868 42424
rect 970 42394 1500 42404
rect 970 42328 980 42394
rect 1490 42328 1500 42394
rect 970 42318 1500 42328
rect 342 42298 868 42308
rect 342 42232 352 42298
rect 858 42232 868 42298
rect 342 42222 868 42232
rect 970 42202 1500 42212
rect 970 42136 980 42202
rect 1490 42136 1500 42202
rect 970 42126 1500 42136
rect 342 42106 868 42116
rect 342 42040 352 42106
rect 858 42040 868 42106
rect 342 42030 868 42040
rect 970 42010 1500 42020
rect 970 41944 980 42010
rect 1490 41944 1500 42010
rect 970 41934 1500 41944
rect 342 41914 868 41924
rect 342 41848 352 41914
rect 858 41848 868 41914
rect 342 41838 868 41848
rect 970 41818 1500 41828
rect 970 41752 980 41818
rect 1490 41752 1500 41818
rect 970 41742 1500 41752
rect 342 41722 868 41732
rect 342 41656 352 41722
rect 858 41656 868 41722
rect 342 41646 868 41656
rect 970 41626 1500 41636
rect 970 41560 980 41626
rect 1490 41560 1500 41626
rect 970 41550 1500 41560
rect 342 41530 868 41540
rect 342 41464 352 41530
rect 858 41464 868 41530
rect 342 41454 868 41464
rect 970 41434 1500 41444
rect 970 41368 980 41434
rect 1490 41368 1500 41434
rect 970 41358 1500 41368
rect 342 41338 868 41348
rect 342 41272 352 41338
rect 858 41272 868 41338
rect 342 41262 868 41272
rect 970 41242 1500 41252
rect 970 41176 980 41242
rect 1490 41176 1500 41242
rect 970 41166 1500 41176
rect 342 41146 868 41156
rect 342 41080 352 41146
rect 858 41080 868 41146
rect 342 41070 868 41080
rect 970 41050 1500 41060
rect 970 40984 980 41050
rect 1490 40984 1500 41050
rect 970 40974 1500 40984
rect 342 40954 868 40964
rect 342 40888 352 40954
rect 858 40888 868 40954
rect 342 40878 868 40888
rect 970 40858 1500 40868
rect 970 40792 980 40858
rect 1490 40792 1500 40858
rect 970 40782 1500 40792
rect 342 40762 868 40772
rect 342 40696 352 40762
rect 858 40696 868 40762
rect 342 40686 868 40696
rect 970 40666 1500 40676
rect 970 40600 980 40666
rect 1490 40600 1500 40666
rect 970 40590 1500 40600
rect 342 40570 868 40580
rect 342 40504 352 40570
rect 858 40504 868 40570
rect 342 40494 868 40504
rect 970 40474 1500 40484
rect 970 40408 980 40474
rect 1490 40408 1500 40474
rect 970 40398 1500 40408
rect 342 40378 868 40388
rect 342 40312 352 40378
rect 858 40312 868 40378
rect 342 40302 868 40312
rect 970 40282 1500 40292
rect 970 40216 980 40282
rect 1490 40216 1500 40282
rect 970 40206 1500 40216
rect 342 40186 868 40196
rect 342 40120 352 40186
rect 858 40120 868 40186
rect 342 40110 868 40120
rect 970 40090 1500 40100
rect 970 40024 980 40090
rect 1490 40024 1500 40090
rect 970 40014 1500 40024
rect 342 39994 868 40004
rect 342 39928 352 39994
rect 858 39928 868 39994
rect 342 39918 868 39928
rect 970 39898 1500 39908
rect 970 39832 980 39898
rect 1490 39832 1500 39898
rect 970 39822 1500 39832
rect 342 39802 868 39812
rect 342 39736 352 39802
rect 858 39736 868 39802
rect 342 39726 868 39736
rect 970 39706 1500 39716
rect 970 39640 980 39706
rect 1490 39640 1500 39706
rect 970 39630 1500 39640
rect 342 39610 868 39620
rect 342 39544 352 39610
rect 858 39544 868 39610
rect 342 39534 868 39544
rect 970 39514 1500 39524
rect 970 39448 980 39514
rect 1490 39448 1500 39514
rect 970 39438 1500 39448
rect 342 39418 868 39428
rect 342 39352 352 39418
rect 858 39352 868 39418
rect 342 39342 868 39352
rect 970 39322 1500 39332
rect 970 39256 980 39322
rect 1490 39256 1500 39322
rect 970 39246 1500 39256
rect 342 39226 868 39236
rect 342 39160 352 39226
rect 858 39160 868 39226
rect 342 39150 868 39160
rect 970 39130 1500 39140
rect 970 39064 980 39130
rect 1490 39064 1500 39130
rect 970 39054 1500 39064
rect 342 39034 868 39044
rect 342 38968 352 39034
rect 858 38968 868 39034
rect 342 38958 868 38968
rect 970 38938 1500 38948
rect 970 38872 980 38938
rect 1490 38872 1500 38938
rect 970 38862 1500 38872
rect 342 38842 868 38852
rect 342 38776 352 38842
rect 858 38776 868 38842
rect 342 38766 868 38776
rect 970 38746 1500 38756
rect 970 38680 980 38746
rect 1490 38680 1500 38746
rect 970 38670 1500 38680
rect 342 38650 868 38660
rect 342 38584 352 38650
rect 858 38584 868 38650
rect 342 38574 868 38584
rect 970 38554 1500 38564
rect 970 38488 980 38554
rect 1490 38488 1500 38554
rect 970 38478 1500 38488
rect 342 38458 868 38468
rect 342 38392 352 38458
rect 858 38392 868 38458
rect 342 38382 868 38392
rect 970 38362 1500 38372
rect 970 38296 980 38362
rect 1490 38296 1500 38362
rect 970 38286 1500 38296
rect 342 38266 868 38276
rect 342 38200 352 38266
rect 858 38200 868 38266
rect 342 38190 868 38200
rect 970 38170 1500 38180
rect 970 38104 980 38170
rect 1490 38104 1500 38170
rect 970 38094 1500 38104
rect 342 38074 868 38084
rect 342 38008 352 38074
rect 858 38008 868 38074
rect 342 37998 868 38008
rect 970 37978 1500 37988
rect 970 37912 980 37978
rect 1490 37912 1500 37978
rect 970 37902 1500 37912
rect 342 37882 868 37892
rect 342 37816 352 37882
rect 858 37816 868 37882
rect 342 37806 868 37816
rect 970 37786 1500 37796
rect 970 37720 980 37786
rect 1490 37720 1500 37786
rect 970 37710 1500 37720
rect 342 37690 868 37700
rect 342 37624 352 37690
rect 858 37624 868 37690
rect 342 37614 868 37624
rect 970 37594 1500 37604
rect 970 37528 980 37594
rect 1490 37528 1500 37594
rect 970 37518 1500 37528
rect 342 37498 868 37508
rect 342 37432 352 37498
rect 858 37432 868 37498
rect 342 37422 868 37432
rect 970 37402 1500 37412
rect 970 37336 980 37402
rect 1490 37336 1500 37402
rect 970 37326 1500 37336
rect 342 37306 868 37316
rect 342 37240 352 37306
rect 858 37240 868 37306
rect 342 37230 868 37240
rect 970 37210 1500 37220
rect 970 37144 980 37210
rect 1490 37144 1500 37210
rect 970 37134 1500 37144
rect 342 37114 868 37124
rect 342 37048 352 37114
rect 858 37048 868 37114
rect 342 37038 868 37048
rect 970 37018 1500 37028
rect 970 36952 980 37018
rect 1490 36952 1500 37018
rect 970 36942 1500 36952
rect 342 36922 868 36932
rect 342 36856 352 36922
rect 858 36856 868 36922
rect 342 36846 868 36856
rect 970 36826 1500 36836
rect 970 36760 980 36826
rect 1490 36760 1500 36826
rect 970 36750 1500 36760
rect 342 36730 868 36740
rect 342 36664 352 36730
rect 858 36664 868 36730
rect 342 36654 868 36664
rect 970 36634 1500 36644
rect 970 36568 980 36634
rect 1490 36568 1500 36634
rect 970 36558 1500 36568
rect 342 36538 868 36548
rect 342 36472 352 36538
rect 858 36472 868 36538
rect 342 36462 868 36472
rect 970 36442 1500 36452
rect 970 36376 980 36442
rect 1490 36376 1500 36442
rect 970 36366 1500 36376
rect 342 36346 868 36356
rect 342 36280 352 36346
rect 858 36280 868 36346
rect 342 36270 868 36280
rect 970 36250 1500 36260
rect 970 36184 980 36250
rect 1490 36184 1500 36250
rect 970 36174 1500 36184
rect 342 36154 868 36164
rect 342 36088 352 36154
rect 858 36088 868 36154
rect 342 36078 868 36088
rect 970 36058 1500 36068
rect 970 35992 980 36058
rect 1490 35992 1500 36058
rect 970 35982 1500 35992
rect 342 35962 868 35972
rect 342 35896 352 35962
rect 858 35896 868 35962
rect 342 35886 868 35896
rect 970 35866 1500 35876
rect 970 35800 980 35866
rect 1490 35800 1500 35866
rect 970 35790 1500 35800
rect 342 35770 868 35780
rect 342 35704 352 35770
rect 858 35704 868 35770
rect 342 35694 868 35704
rect 970 35674 1500 35684
rect 970 35608 980 35674
rect 1490 35608 1500 35674
rect 970 35598 1500 35608
rect 342 35578 868 35588
rect 342 35512 352 35578
rect 858 35512 868 35578
rect 342 35502 868 35512
rect 970 35482 1500 35492
rect 970 35416 980 35482
rect 1490 35416 1500 35482
rect 970 35406 1500 35416
rect 342 35386 868 35396
rect 342 35320 352 35386
rect 858 35320 868 35386
rect 342 35310 868 35320
rect 970 35290 1500 35300
rect 970 35224 980 35290
rect 1490 35224 1500 35290
rect 970 35214 1500 35224
rect 342 35194 868 35204
rect 342 35128 352 35194
rect 858 35128 868 35194
rect 342 35118 868 35128
rect 970 35098 1500 35108
rect 970 35032 980 35098
rect 1490 35032 1500 35098
rect 970 35022 1500 35032
rect 342 35002 868 35012
rect 342 34936 352 35002
rect 858 34936 868 35002
rect 342 34926 868 34936
rect 970 34906 1500 34916
rect 970 34840 980 34906
rect 1490 34840 1500 34906
rect 970 34830 1500 34840
rect 342 34810 868 34820
rect 342 34744 352 34810
rect 858 34744 868 34810
rect 342 34734 868 34744
rect 970 34714 1500 34724
rect 970 34648 980 34714
rect 1490 34648 1500 34714
rect 970 34638 1500 34648
rect 342 34618 868 34628
rect 342 34552 352 34618
rect 858 34552 868 34618
rect 342 34542 868 34552
rect 970 34522 1500 34532
rect 970 34456 980 34522
rect 1490 34456 1500 34522
rect 970 34446 1500 34456
rect 342 34426 868 34436
rect 342 34360 352 34426
rect 858 34360 868 34426
rect 342 34350 868 34360
rect 970 34330 1500 34340
rect 970 34264 980 34330
rect 1490 34264 1500 34330
rect 970 34254 1500 34264
rect 342 34234 868 34244
rect 342 34168 352 34234
rect 858 34168 868 34234
rect 342 34158 868 34168
rect 970 34138 1500 34148
rect 970 34072 980 34138
rect 1490 34072 1500 34138
rect 970 34062 1500 34072
rect 342 34042 868 34052
rect 342 33976 352 34042
rect 858 33976 868 34042
rect 342 33966 868 33976
rect 970 33946 1500 33956
rect 970 33880 980 33946
rect 1490 33880 1500 33946
rect 970 33870 1500 33880
rect 342 33850 868 33860
rect 342 33784 352 33850
rect 858 33784 868 33850
rect 342 33774 868 33784
rect 970 33754 1500 33764
rect 970 33688 980 33754
rect 1490 33688 1500 33754
rect 970 33678 1500 33688
rect 342 33658 868 33668
rect 342 33592 352 33658
rect 858 33592 868 33658
rect 342 33582 868 33592
rect 970 33562 1500 33572
rect 970 33496 980 33562
rect 1490 33496 1500 33562
rect 970 33486 1500 33496
rect 342 33466 868 33476
rect 342 33400 352 33466
rect 858 33400 868 33466
rect 342 33390 868 33400
rect 970 33370 1500 33380
rect 970 33304 980 33370
rect 1490 33304 1500 33370
rect 970 33294 1500 33304
rect 342 33274 868 33284
rect 342 33208 352 33274
rect 858 33208 868 33274
rect 342 33198 868 33208
rect 970 33178 1500 33188
rect 970 33112 980 33178
rect 1490 33112 1500 33178
rect 970 33102 1500 33112
rect 342 33082 868 33092
rect 342 33016 352 33082
rect 858 33016 868 33082
rect 342 33006 868 33016
rect 970 32986 1500 32996
rect 970 32920 980 32986
rect 1490 32920 1500 32986
rect 970 32910 1500 32920
rect 342 32890 868 32900
rect 342 32824 352 32890
rect 858 32824 868 32890
rect 342 32814 868 32824
rect 970 32794 1500 32804
rect 970 32728 980 32794
rect 1490 32728 1500 32794
rect 970 32718 1500 32728
rect 342 32698 868 32708
rect 342 32632 352 32698
rect 858 32632 868 32698
rect 342 32622 868 32632
rect 970 32602 1500 32612
rect 970 32536 980 32602
rect 1490 32536 1500 32602
rect 970 32526 1500 32536
rect 342 32506 868 32516
rect 342 32440 352 32506
rect 858 32440 868 32506
rect 342 32430 868 32440
rect 970 32410 1500 32420
rect 970 32344 980 32410
rect 1490 32344 1500 32410
rect 970 32334 1500 32344
rect 342 32314 868 32324
rect 342 32248 352 32314
rect 858 32248 868 32314
rect 342 32238 868 32248
rect 970 32218 1500 32228
rect 970 32152 980 32218
rect 1490 32152 1500 32218
rect 970 32142 1500 32152
rect 342 32122 868 32132
rect 342 32056 352 32122
rect 858 32056 868 32122
rect 342 32046 868 32056
rect 970 32026 1500 32036
rect 970 31960 980 32026
rect 1490 31960 1500 32026
rect 970 31950 1500 31960
rect 342 31930 868 31940
rect 342 31864 352 31930
rect 858 31864 868 31930
rect 342 31854 868 31864
rect 970 31834 1500 31844
rect 970 31768 980 31834
rect 1490 31768 1500 31834
rect 970 31758 1500 31768
rect 342 31738 868 31748
rect 342 31672 352 31738
rect 858 31672 868 31738
rect 342 31662 868 31672
rect 970 31642 1500 31652
rect 970 31576 980 31642
rect 1490 31576 1500 31642
rect 970 31566 1500 31576
rect 342 31546 868 31556
rect 342 31480 352 31546
rect 858 31480 868 31546
rect 342 31470 868 31480
rect 970 31450 1500 31460
rect 970 31384 980 31450
rect 1490 31384 1500 31450
rect 970 31374 1500 31384
rect 342 31354 868 31364
rect 342 31288 352 31354
rect 858 31288 868 31354
rect 342 31278 868 31288
rect 970 31258 1500 31268
rect 970 31192 980 31258
rect 1490 31192 1500 31258
rect 970 31182 1500 31192
rect 342 31162 868 31172
rect 342 31096 352 31162
rect 858 31096 868 31162
rect 342 31086 868 31096
rect 970 31066 1500 31076
rect 970 31000 980 31066
rect 1490 31000 1500 31066
rect 970 30990 1500 31000
rect 342 30970 868 30980
rect 342 30904 352 30970
rect 858 30904 868 30970
rect 342 30894 868 30904
rect 970 30874 1500 30884
rect 970 30808 980 30874
rect 1490 30808 1500 30874
rect 970 30798 1500 30808
rect 342 30778 868 30788
rect 342 30712 352 30778
rect 858 30712 868 30778
rect 342 30702 868 30712
rect 970 30682 1500 30692
rect 970 30616 980 30682
rect 1490 30616 1500 30682
rect 970 30606 1500 30616
rect 342 30586 868 30596
rect 342 30520 352 30586
rect 858 30520 868 30586
rect 342 30510 868 30520
rect 970 30490 1500 30500
rect 970 30424 980 30490
rect 1490 30424 1500 30490
rect 970 30414 1500 30424
rect 342 30394 868 30404
rect 342 30328 352 30394
rect 858 30328 868 30394
rect 342 30318 868 30328
rect 970 30298 1500 30308
rect 970 30232 980 30298
rect 1490 30232 1500 30298
rect 970 30222 1500 30232
rect 342 30202 868 30212
rect 342 30136 352 30202
rect 858 30136 868 30202
rect 342 30126 868 30136
rect 970 30106 1500 30116
rect 970 30040 980 30106
rect 1490 30040 1500 30106
rect 970 30030 1500 30040
rect 342 30010 868 30020
rect 342 29944 352 30010
rect 858 29944 868 30010
rect 342 29934 868 29944
rect 970 29914 1500 29924
rect 970 29848 980 29914
rect 1490 29848 1500 29914
rect 970 29838 1500 29848
rect 342 29818 868 29828
rect 342 29752 352 29818
rect 858 29752 868 29818
rect 342 29742 868 29752
rect 970 29722 1500 29732
rect 970 29656 980 29722
rect 1490 29656 1500 29722
rect 970 29646 1500 29656
rect 342 29626 868 29636
rect 342 29560 352 29626
rect 858 29560 868 29626
rect 342 29550 868 29560
rect 970 29530 1500 29540
rect 970 29464 980 29530
rect 1490 29464 1500 29530
rect 970 29454 1500 29464
rect 342 29434 868 29444
rect 342 29368 352 29434
rect 858 29368 868 29434
rect 342 29358 868 29368
rect 970 29338 1500 29348
rect 970 29272 980 29338
rect 1490 29272 1500 29338
rect 970 29262 1500 29272
rect 342 29242 868 29252
rect 342 29176 352 29242
rect 858 29176 868 29242
rect 342 29166 868 29176
rect 970 29146 1500 29156
rect 970 29080 980 29146
rect 1490 29080 1500 29146
rect 970 29070 1500 29080
rect 342 29050 868 29060
rect 342 28984 352 29050
rect 858 28984 868 29050
rect 342 28974 868 28984
rect 970 28954 1500 28964
rect 970 28888 980 28954
rect 1490 28888 1500 28954
rect 970 28878 1500 28888
rect 342 28858 868 28868
rect 342 28792 352 28858
rect 858 28792 868 28858
rect 342 28782 868 28792
rect 970 28762 1500 28772
rect 970 28696 980 28762
rect 1490 28696 1500 28762
rect 970 28686 1500 28696
rect 342 28666 868 28676
rect 342 28600 352 28666
rect 858 28600 868 28666
rect 342 28590 868 28600
rect 970 28570 1500 28580
rect 970 28504 980 28570
rect 1490 28504 1500 28570
rect 970 28494 1500 28504
rect 342 28474 868 28484
rect 342 28408 352 28474
rect 858 28408 868 28474
rect 342 28398 868 28408
rect 970 28378 1500 28388
rect 970 28312 980 28378
rect 1490 28312 1500 28378
rect 970 28302 1500 28312
rect 342 28282 868 28292
rect 342 28216 352 28282
rect 858 28216 868 28282
rect 342 28206 868 28216
rect 970 28186 1500 28196
rect 970 28120 980 28186
rect 1490 28120 1500 28186
rect 970 28110 1500 28120
rect 342 28090 868 28100
rect 342 28024 352 28090
rect 858 28024 868 28090
rect 342 28014 868 28024
rect 970 27994 1500 28004
rect 970 27928 980 27994
rect 1490 27928 1500 27994
rect 970 27918 1500 27928
rect 342 27898 868 27908
rect 342 27832 352 27898
rect 858 27832 868 27898
rect 342 27822 868 27832
rect 970 27802 1500 27812
rect 970 27736 980 27802
rect 1490 27736 1500 27802
rect 970 27726 1500 27736
rect 342 27706 868 27716
rect 342 27640 352 27706
rect 858 27640 868 27706
rect 342 27630 868 27640
rect 970 27610 1500 27620
rect 970 27544 980 27610
rect 1490 27544 1500 27610
rect 970 27534 1500 27544
rect 342 27514 868 27524
rect 342 27448 352 27514
rect 858 27448 868 27514
rect 342 27438 868 27448
rect 970 27418 1500 27428
rect 970 27352 980 27418
rect 1490 27352 1500 27418
rect 970 27342 1500 27352
rect 342 27322 868 27332
rect 342 27256 352 27322
rect 858 27256 868 27322
rect 342 27246 868 27256
rect 970 27226 1500 27236
rect 970 27160 980 27226
rect 1490 27160 1500 27226
rect 970 27150 1500 27160
rect 342 27130 868 27140
rect 342 27064 352 27130
rect 858 27064 868 27130
rect 342 27054 868 27064
rect 970 27034 1500 27044
rect 970 26968 980 27034
rect 1490 26968 1500 27034
rect 970 26958 1500 26968
rect 342 26938 868 26948
rect 342 26872 352 26938
rect 858 26872 868 26938
rect 342 26862 868 26872
rect 970 26842 1500 26852
rect 970 26776 980 26842
rect 1490 26776 1500 26842
rect 970 26766 1500 26776
rect 342 26746 868 26756
rect 342 26680 352 26746
rect 858 26680 868 26746
rect 342 26670 868 26680
rect 970 26650 1500 26660
rect 970 26584 980 26650
rect 1490 26584 1500 26650
rect 970 26574 1500 26584
rect 342 26554 868 26564
rect 342 26488 352 26554
rect 858 26488 868 26554
rect 342 26478 868 26488
rect 970 26458 1500 26468
rect 970 26392 980 26458
rect 1490 26392 1500 26458
rect 970 26382 1500 26392
rect 342 26362 868 26372
rect 342 26296 352 26362
rect 858 26296 868 26362
rect 342 26286 868 26296
rect 970 26266 1500 26276
rect 970 26200 980 26266
rect 1490 26200 1500 26266
rect 970 26190 1500 26200
rect 342 26170 868 26180
rect 342 26104 352 26170
rect 858 26104 868 26170
rect 342 26094 868 26104
rect 970 26074 1500 26084
rect 970 26008 980 26074
rect 1490 26008 1500 26074
rect 970 25998 1500 26008
rect 342 25978 868 25988
rect 342 25912 352 25978
rect 858 25912 868 25978
rect 342 25902 868 25912
rect 970 25882 1500 25892
rect 970 25816 980 25882
rect 1490 25816 1500 25882
rect 970 25806 1500 25816
rect 342 25786 868 25796
rect 342 25720 352 25786
rect 858 25720 868 25786
rect 342 25710 868 25720
rect 970 25690 1500 25700
rect 970 25624 980 25690
rect 1490 25624 1500 25690
rect 970 25614 1500 25624
rect 342 25594 868 25604
rect 342 25528 352 25594
rect 858 25528 868 25594
rect 342 25518 868 25528
rect 970 25498 1500 25508
rect 970 25432 980 25498
rect 1490 25432 1500 25498
rect 970 25422 1500 25432
rect 342 25402 868 25412
rect 342 25336 352 25402
rect 858 25336 868 25402
rect 342 25326 868 25336
rect 970 25306 1500 25316
rect 970 25240 980 25306
rect 1490 25240 1500 25306
rect 970 25230 1500 25240
rect 342 25210 868 25220
rect 342 25144 352 25210
rect 858 25144 868 25210
rect 342 25134 868 25144
rect 970 25114 1500 25124
rect 970 25048 980 25114
rect 1490 25048 1500 25114
rect 970 25038 1500 25048
rect 342 25018 868 25028
rect 342 24952 352 25018
rect 858 24952 868 25018
rect 342 24942 868 24952
rect 970 24922 1500 24932
rect 970 24856 980 24922
rect 1490 24856 1500 24922
rect 970 24846 1500 24856
rect 342 24826 868 24836
rect 342 24760 352 24826
rect 858 24760 868 24826
rect 342 24750 868 24760
rect 970 24730 1500 24740
rect 970 24664 980 24730
rect 1490 24664 1500 24730
rect 970 24654 1500 24664
rect 342 24634 868 24644
rect 342 24568 352 24634
rect 858 24568 868 24634
rect 342 24558 868 24568
rect 970 24538 1500 24548
rect 970 24472 980 24538
rect 1490 24472 1500 24538
rect 970 24462 1500 24472
rect 342 24442 868 24452
rect 342 24376 352 24442
rect 858 24376 868 24442
rect 342 24366 868 24376
rect 970 24346 1500 24356
rect 970 24280 980 24346
rect 1490 24280 1500 24346
rect 970 24270 1500 24280
rect 342 24250 868 24260
rect 342 24184 352 24250
rect 858 24184 868 24250
rect 342 24174 868 24184
rect 970 24154 1500 24164
rect 970 24088 980 24154
rect 1490 24088 1500 24154
rect 970 24078 1500 24088
rect 342 24058 868 24068
rect 342 23992 352 24058
rect 858 23992 868 24058
rect 342 23982 868 23992
rect 970 23962 1500 23972
rect 970 23896 980 23962
rect 1490 23896 1500 23962
rect 970 23886 1500 23896
rect 342 23866 868 23876
rect 342 23800 352 23866
rect 858 23800 868 23866
rect 342 23790 868 23800
rect 970 23770 1500 23780
rect 970 23704 980 23770
rect 1490 23704 1500 23770
rect 970 23694 1500 23704
rect 342 23674 868 23684
rect 342 23608 352 23674
rect 858 23608 868 23674
rect 342 23598 868 23608
rect 970 23578 1500 23588
rect 970 23512 980 23578
rect 1490 23512 1500 23578
rect 970 23502 1500 23512
rect 342 23482 868 23492
rect 342 23416 352 23482
rect 858 23416 868 23482
rect 342 23406 868 23416
rect 970 23386 1500 23396
rect 970 23320 980 23386
rect 1490 23320 1500 23386
rect 970 23310 1500 23320
rect 342 23290 868 23300
rect 342 23224 352 23290
rect 858 23224 868 23290
rect 342 23214 868 23224
rect 970 23194 1500 23204
rect 970 23128 980 23194
rect 1490 23128 1500 23194
rect 970 23118 1500 23128
rect 342 23098 868 23108
rect 342 23032 352 23098
rect 858 23032 868 23098
rect 342 23022 868 23032
rect 330 22768 880 22773
rect 330 21986 340 22768
rect 870 21986 880 22768
rect 330 21981 880 21986
rect 342 21720 868 21730
rect 342 21654 352 21720
rect 858 21654 868 21720
rect 342 21644 868 21654
rect 970 21624 1500 21634
rect 970 21558 980 21624
rect 1490 21558 1500 21624
rect 970 21548 1500 21558
rect 342 21528 868 21538
rect 342 21462 352 21528
rect 858 21462 868 21528
rect 342 21452 868 21462
rect 970 21432 1500 21442
rect 970 21366 980 21432
rect 1490 21366 1500 21432
rect 970 21356 1500 21366
rect 342 21336 868 21346
rect 342 21270 352 21336
rect 858 21270 868 21336
rect 342 21260 868 21270
rect 970 21240 1500 21250
rect 970 21174 980 21240
rect 1490 21174 1500 21240
rect 970 21164 1500 21174
rect 342 21144 868 21154
rect 342 21078 352 21144
rect 858 21078 868 21144
rect 342 21068 868 21078
rect 970 21048 1500 21058
rect 970 20982 980 21048
rect 1490 20982 1500 21048
rect 970 20972 1500 20982
rect 342 20952 868 20962
rect 342 20886 352 20952
rect 858 20886 868 20952
rect 342 20876 868 20886
rect 970 20856 1500 20866
rect 970 20790 980 20856
rect 1490 20790 1500 20856
rect 970 20780 1500 20790
rect 342 20760 868 20770
rect 342 20694 352 20760
rect 858 20694 868 20760
rect 342 20684 868 20694
rect 970 20664 1500 20674
rect 970 20598 980 20664
rect 1490 20598 1500 20664
rect 970 20588 1500 20598
rect 342 20568 868 20578
rect 342 20502 352 20568
rect 858 20502 868 20568
rect 342 20492 868 20502
rect 970 20472 1500 20482
rect 970 20406 980 20472
rect 1490 20406 1500 20472
rect 970 20396 1500 20406
rect 342 20376 868 20386
rect 342 20310 352 20376
rect 858 20310 868 20376
rect 342 20300 868 20310
rect 970 20280 1500 20290
rect 970 20214 980 20280
rect 1490 20214 1500 20280
rect 970 20204 1500 20214
rect 342 20184 868 20194
rect 342 20118 352 20184
rect 858 20118 868 20184
rect 342 20108 868 20118
rect 970 20088 1500 20098
rect 970 20022 980 20088
rect 1490 20022 1500 20088
rect 970 20012 1500 20022
rect 342 19992 868 20002
rect 342 19926 352 19992
rect 858 19926 868 19992
rect 342 19916 868 19926
rect 970 19896 1500 19906
rect 970 19830 980 19896
rect 1490 19830 1500 19896
rect 970 19820 1500 19830
rect 342 19800 868 19810
rect 342 19734 352 19800
rect 858 19734 868 19800
rect 342 19724 868 19734
rect 970 19704 1500 19714
rect 970 19638 980 19704
rect 1490 19638 1500 19704
rect 970 19628 1500 19638
rect 342 19608 868 19618
rect 342 19542 352 19608
rect 858 19542 868 19608
rect 342 19532 868 19542
rect 970 19512 1500 19522
rect 970 19446 980 19512
rect 1490 19446 1500 19512
rect 970 19436 1500 19446
rect 342 19416 868 19426
rect 342 19350 352 19416
rect 858 19350 868 19416
rect 342 19340 868 19350
rect 970 19320 1500 19330
rect 970 19254 980 19320
rect 1490 19254 1500 19320
rect 970 19244 1500 19254
rect 342 19224 868 19234
rect 342 19158 352 19224
rect 858 19158 868 19224
rect 342 19148 868 19158
rect 970 19128 1500 19138
rect 970 19062 980 19128
rect 1490 19062 1500 19128
rect 970 19052 1500 19062
rect 342 19032 868 19042
rect 342 18966 352 19032
rect 858 18966 868 19032
rect 342 18956 868 18966
rect 970 18936 1500 18946
rect 970 18870 980 18936
rect 1490 18870 1500 18936
rect 970 18860 1500 18870
rect 342 18840 868 18850
rect 342 18774 352 18840
rect 858 18774 868 18840
rect 342 18764 868 18774
rect 970 18744 1500 18754
rect 970 18678 980 18744
rect 1490 18678 1500 18744
rect 970 18668 1500 18678
rect 342 18648 868 18658
rect 342 18582 352 18648
rect 858 18582 868 18648
rect 342 18572 868 18582
rect 970 18552 1500 18562
rect 970 18486 980 18552
rect 1490 18486 1500 18552
rect 970 18476 1500 18486
rect 342 18456 868 18466
rect 342 18390 352 18456
rect 858 18390 868 18456
rect 342 18380 868 18390
rect 970 18360 1500 18370
rect 970 18294 980 18360
rect 1490 18294 1500 18360
rect 970 18284 1500 18294
rect 342 18264 868 18274
rect 342 18198 352 18264
rect 858 18198 868 18264
rect 342 18188 868 18198
rect 970 18168 1500 18178
rect 970 18102 980 18168
rect 1490 18102 1500 18168
rect 970 18092 1500 18102
rect 342 18072 868 18082
rect 342 18006 352 18072
rect 858 18006 868 18072
rect 342 17996 868 18006
rect 970 17976 1500 17986
rect 970 17910 980 17976
rect 1490 17910 1500 17976
rect 970 17900 1500 17910
rect 342 17880 868 17890
rect 342 17814 352 17880
rect 858 17814 868 17880
rect 342 17804 868 17814
rect 970 17784 1500 17794
rect 970 17718 980 17784
rect 1490 17718 1500 17784
rect 970 17708 1500 17718
rect 342 17688 868 17698
rect 342 17622 352 17688
rect 858 17622 868 17688
rect 342 17612 868 17622
rect 970 17592 1500 17602
rect 970 17526 980 17592
rect 1490 17526 1500 17592
rect 970 17516 1500 17526
rect 342 17496 868 17506
rect 342 17430 352 17496
rect 858 17430 868 17496
rect 342 17420 868 17430
rect 970 17400 1500 17410
rect 970 17334 980 17400
rect 1490 17334 1500 17400
rect 970 17324 1500 17334
rect 342 17304 868 17314
rect 342 17238 352 17304
rect 858 17238 868 17304
rect 342 17228 868 17238
rect 970 17208 1500 17218
rect 970 17142 980 17208
rect 1490 17142 1500 17208
rect 970 17132 1500 17142
rect 342 17112 868 17122
rect 342 17046 352 17112
rect 858 17046 868 17112
rect 342 17036 868 17046
rect 970 17016 1500 17026
rect 970 16950 980 17016
rect 1490 16950 1500 17016
rect 970 16940 1500 16950
rect 342 16920 868 16930
rect 342 16854 352 16920
rect 858 16854 868 16920
rect 342 16844 868 16854
rect 970 16824 1500 16834
rect 970 16758 980 16824
rect 1490 16758 1500 16824
rect 970 16748 1500 16758
rect 342 16728 868 16738
rect 342 16662 352 16728
rect 858 16662 868 16728
rect 342 16652 868 16662
rect 970 16632 1500 16642
rect 970 16566 980 16632
rect 1490 16566 1500 16632
rect 970 16556 1500 16566
rect 342 16536 868 16546
rect 342 16470 352 16536
rect 858 16470 868 16536
rect 342 16460 868 16470
rect 970 16440 1500 16450
rect 970 16374 980 16440
rect 1490 16374 1500 16440
rect 970 16364 1500 16374
rect 342 16344 868 16354
rect 342 16278 352 16344
rect 858 16278 868 16344
rect 342 16268 868 16278
rect 970 16248 1500 16258
rect 970 16182 980 16248
rect 1490 16182 1500 16248
rect 970 16172 1500 16182
rect 342 16152 868 16162
rect 342 16086 352 16152
rect 858 16086 868 16152
rect 342 16076 868 16086
rect 970 16056 1500 16066
rect 970 15990 980 16056
rect 1490 15990 1500 16056
rect 970 15980 1500 15990
rect 342 15960 868 15970
rect 342 15894 352 15960
rect 858 15894 868 15960
rect 342 15884 868 15894
rect 970 15864 1500 15874
rect 970 15798 980 15864
rect 1490 15798 1500 15864
rect 970 15788 1500 15798
rect 342 15768 868 15778
rect 342 15702 352 15768
rect 858 15702 868 15768
rect 342 15692 868 15702
rect 970 15672 1500 15682
rect 970 15606 980 15672
rect 1490 15606 1500 15672
rect 970 15596 1500 15606
rect 342 15576 868 15586
rect 342 15510 352 15576
rect 858 15510 868 15576
rect 342 15500 868 15510
rect 970 15480 1500 15490
rect 970 15414 980 15480
rect 1490 15414 1500 15480
rect 970 15404 1500 15414
rect 342 15384 868 15394
rect 342 15318 352 15384
rect 858 15318 868 15384
rect 342 15308 868 15318
rect 970 15288 1500 15298
rect 970 15222 980 15288
rect 1490 15222 1500 15288
rect 970 15212 1500 15222
rect 342 15192 868 15202
rect 342 15126 352 15192
rect 858 15126 868 15192
rect 342 15116 868 15126
rect 970 15096 1500 15106
rect 970 15030 980 15096
rect 1490 15030 1500 15096
rect 970 15020 1500 15030
rect 342 15000 868 15010
rect 342 14934 352 15000
rect 858 14934 868 15000
rect 342 14924 868 14934
rect 970 14904 1500 14914
rect 970 14838 980 14904
rect 1490 14838 1500 14904
rect 970 14828 1500 14838
rect 342 14808 868 14818
rect 342 14742 352 14808
rect 858 14742 868 14808
rect 342 14732 868 14742
rect 970 14712 1500 14722
rect 970 14646 980 14712
rect 1490 14646 1500 14712
rect 970 14636 1500 14646
rect 342 14616 868 14626
rect 342 14550 352 14616
rect 858 14550 868 14616
rect 342 14540 868 14550
rect 970 14520 1500 14530
rect 970 14454 980 14520
rect 1490 14454 1500 14520
rect 970 14444 1500 14454
rect 342 14424 868 14434
rect 342 14358 352 14424
rect 858 14358 868 14424
rect 342 14348 868 14358
rect 970 14328 1500 14338
rect 970 14262 980 14328
rect 1490 14262 1500 14328
rect 970 14252 1500 14262
rect 342 14232 868 14242
rect 342 14166 352 14232
rect 858 14166 868 14232
rect 342 14156 868 14166
rect 970 14136 1500 14146
rect 970 14070 980 14136
rect 1490 14070 1500 14136
rect 970 14060 1500 14070
rect 342 14040 868 14050
rect 342 13974 352 14040
rect 858 13974 868 14040
rect 342 13964 868 13974
rect 970 13944 1500 13954
rect 970 13878 980 13944
rect 1490 13878 1500 13944
rect 970 13868 1500 13878
rect 342 13848 868 13858
rect 342 13782 352 13848
rect 858 13782 868 13848
rect 342 13772 868 13782
rect 970 13752 1500 13762
rect 970 13686 980 13752
rect 1490 13686 1500 13752
rect 970 13676 1500 13686
rect 342 13656 868 13666
rect 342 13590 352 13656
rect 858 13590 868 13656
rect 342 13580 868 13590
rect 970 13560 1500 13570
rect 970 13494 980 13560
rect 1490 13494 1500 13560
rect 970 13484 1500 13494
rect 342 13464 868 13474
rect 342 13398 352 13464
rect 858 13398 868 13464
rect 342 13388 868 13398
rect 970 13368 1500 13378
rect 970 13302 980 13368
rect 1490 13302 1500 13368
rect 970 13292 1500 13302
rect 342 13272 868 13282
rect 342 13206 352 13272
rect 858 13206 868 13272
rect 342 13196 868 13206
rect 970 13176 1500 13186
rect 970 13110 980 13176
rect 1490 13110 1500 13176
rect 970 13100 1500 13110
rect 342 13080 868 13090
rect 342 13014 352 13080
rect 858 13014 868 13080
rect 342 13004 868 13014
rect 970 12984 1500 12994
rect 970 12918 980 12984
rect 1490 12918 1500 12984
rect 970 12908 1500 12918
rect 342 12888 868 12898
rect 342 12822 352 12888
rect 858 12822 868 12888
rect 342 12812 868 12822
rect 970 12792 1500 12802
rect 970 12726 980 12792
rect 1490 12726 1500 12792
rect 970 12716 1500 12726
rect 342 12696 868 12706
rect 342 12630 352 12696
rect 858 12630 868 12696
rect 342 12620 868 12630
rect 970 12600 1500 12610
rect 970 12534 980 12600
rect 1490 12534 1500 12600
rect 970 12524 1500 12534
rect 342 12504 868 12514
rect 342 12438 352 12504
rect 858 12438 868 12504
rect 342 12428 868 12438
rect 970 12408 1500 12418
rect 970 12342 980 12408
rect 1490 12342 1500 12408
rect 970 12332 1500 12342
rect 342 12312 868 12322
rect 342 12246 352 12312
rect 858 12246 868 12312
rect 342 12236 868 12246
rect 970 12216 1500 12226
rect 970 12150 980 12216
rect 1490 12150 1500 12216
rect 970 12140 1500 12150
rect 342 12120 868 12130
rect 342 12054 352 12120
rect 858 12054 868 12120
rect 342 12044 868 12054
rect 970 12024 1500 12034
rect 970 11958 980 12024
rect 1490 11958 1500 12024
rect 970 11948 1500 11958
rect 342 11928 868 11938
rect 342 11862 352 11928
rect 858 11862 868 11928
rect 342 11852 868 11862
rect 970 11832 1500 11842
rect 970 11766 980 11832
rect 1490 11766 1500 11832
rect 970 11756 1500 11766
rect 342 11736 868 11746
rect 342 11670 352 11736
rect 858 11670 868 11736
rect 342 11660 868 11670
rect 970 11640 1500 11650
rect 970 11574 980 11640
rect 1490 11574 1500 11640
rect 970 11564 1500 11574
rect 342 11544 868 11554
rect 342 11478 352 11544
rect 858 11478 868 11544
rect 342 11468 868 11478
rect 970 11448 1500 11458
rect 970 11382 980 11448
rect 1490 11382 1500 11448
rect 970 11372 1500 11382
rect 342 11352 868 11362
rect 342 11286 352 11352
rect 858 11286 868 11352
rect 342 11276 868 11286
rect 970 11256 1500 11266
rect 970 11190 980 11256
rect 1490 11190 1500 11256
rect 970 11180 1500 11190
rect 342 11160 868 11170
rect 342 11094 352 11160
rect 858 11094 868 11160
rect 342 11084 868 11094
rect 970 11064 1500 11074
rect 970 10998 980 11064
rect 1490 10998 1500 11064
rect 970 10988 1500 10998
rect 342 10968 868 10978
rect 342 10902 352 10968
rect 858 10902 868 10968
rect 342 10892 868 10902
rect 970 10872 1500 10882
rect 970 10806 980 10872
rect 1490 10806 1500 10872
rect 970 10796 1500 10806
rect 342 10776 868 10786
rect 342 10710 352 10776
rect 858 10710 868 10776
rect 342 10700 868 10710
rect 970 10680 1500 10690
rect 970 10614 980 10680
rect 1490 10614 1500 10680
rect 970 10604 1500 10614
rect 342 10584 868 10594
rect 342 10518 352 10584
rect 858 10518 868 10584
rect 342 10508 868 10518
rect 970 10488 1500 10498
rect 970 10422 980 10488
rect 1490 10422 1500 10488
rect 970 10412 1500 10422
rect 342 10392 868 10402
rect 342 10326 352 10392
rect 858 10326 868 10392
rect 342 10316 868 10326
rect 970 10296 1500 10306
rect 970 10230 980 10296
rect 1490 10230 1500 10296
rect 970 10220 1500 10230
rect 342 10200 868 10210
rect 342 10134 352 10200
rect 858 10134 868 10200
rect 342 10124 868 10134
rect 970 10104 1500 10114
rect 970 10038 980 10104
rect 1490 10038 1500 10104
rect 970 10028 1500 10038
rect 342 10008 868 10018
rect 342 9942 352 10008
rect 858 9942 868 10008
rect 342 9932 868 9942
rect 970 9912 1500 9922
rect 970 9846 980 9912
rect 1490 9846 1500 9912
rect 970 9836 1500 9846
rect 342 9816 868 9826
rect 342 9750 352 9816
rect 858 9750 868 9816
rect 342 9740 868 9750
rect 970 9720 1500 9730
rect 970 9654 980 9720
rect 1490 9654 1500 9720
rect 970 9644 1500 9654
rect 342 9624 868 9634
rect 342 9558 352 9624
rect 858 9558 868 9624
rect 342 9548 868 9558
rect 970 9528 1500 9538
rect 970 9462 980 9528
rect 1490 9462 1500 9528
rect 970 9452 1500 9462
rect 342 9432 868 9442
rect 342 9366 352 9432
rect 858 9366 868 9432
rect 342 9356 868 9366
rect 970 9336 1500 9346
rect 970 9270 980 9336
rect 1490 9270 1500 9336
rect 970 9260 1500 9270
rect 342 9240 868 9250
rect 342 9174 352 9240
rect 858 9174 868 9240
rect 342 9164 868 9174
rect 970 9144 1500 9154
rect 970 9078 980 9144
rect 1490 9078 1500 9144
rect 970 9068 1500 9078
rect 342 9048 868 9058
rect 342 8982 352 9048
rect 858 8982 868 9048
rect 342 8972 868 8982
rect 970 8952 1500 8962
rect 970 8886 980 8952
rect 1490 8886 1500 8952
rect 970 8876 1500 8886
rect 342 8856 868 8866
rect 342 8790 352 8856
rect 858 8790 868 8856
rect 342 8780 868 8790
rect 970 8760 1500 8770
rect 970 8694 980 8760
rect 1490 8694 1500 8760
rect 970 8684 1500 8694
rect 342 8664 868 8674
rect 342 8598 352 8664
rect 858 8598 868 8664
rect 342 8588 868 8598
rect 970 8568 1500 8578
rect 970 8502 980 8568
rect 1490 8502 1500 8568
rect 970 8492 1500 8502
rect 342 8472 868 8482
rect 342 8406 352 8472
rect 858 8406 868 8472
rect 342 8396 868 8406
rect 970 8376 1500 8386
rect 970 8310 980 8376
rect 1490 8310 1500 8376
rect 970 8300 1500 8310
rect 342 8280 868 8290
rect 342 8214 352 8280
rect 858 8214 868 8280
rect 342 8204 868 8214
rect 970 8184 1500 8194
rect 970 8118 980 8184
rect 1490 8118 1500 8184
rect 970 8108 1500 8118
rect 342 8088 868 8098
rect 342 8022 352 8088
rect 858 8022 868 8088
rect 342 8012 868 8022
rect 970 7992 1500 8002
rect 970 7926 980 7992
rect 1490 7926 1500 7992
rect 970 7916 1500 7926
rect 342 7896 868 7906
rect 342 7830 352 7896
rect 858 7830 868 7896
rect 342 7820 868 7830
rect 970 7800 1500 7810
rect 970 7734 980 7800
rect 1490 7734 1500 7800
rect 970 7724 1500 7734
rect 342 7704 868 7714
rect 342 7638 352 7704
rect 858 7638 868 7704
rect 342 7628 868 7638
rect 970 7608 1500 7618
rect 970 7542 980 7608
rect 1490 7542 1500 7608
rect 970 7532 1500 7542
rect 342 7512 868 7522
rect 342 7446 352 7512
rect 858 7446 868 7512
rect 342 7436 868 7446
rect 970 7416 1500 7426
rect 970 7350 980 7416
rect 1490 7350 1500 7416
rect 970 7340 1500 7350
rect 342 7320 868 7330
rect 342 7254 352 7320
rect 858 7254 868 7320
rect 342 7244 868 7254
rect 970 7224 1500 7234
rect 970 7158 980 7224
rect 1490 7158 1500 7224
rect 970 7148 1500 7158
rect 342 7128 868 7138
rect 342 7062 352 7128
rect 858 7062 868 7128
rect 342 7052 868 7062
rect 970 7032 1500 7042
rect 970 6966 980 7032
rect 1490 6966 1500 7032
rect 970 6956 1500 6966
rect 342 6936 868 6946
rect 342 6870 352 6936
rect 858 6870 868 6936
rect 342 6860 868 6870
rect 970 6840 1500 6850
rect 970 6774 980 6840
rect 1490 6774 1500 6840
rect 970 6764 1500 6774
rect 342 6744 868 6754
rect 342 6678 352 6744
rect 858 6678 868 6744
rect 342 6668 868 6678
rect 970 6648 1500 6658
rect 970 6582 980 6648
rect 1490 6582 1500 6648
rect 970 6572 1500 6582
rect 342 6552 868 6562
rect 342 6486 352 6552
rect 858 6486 868 6552
rect 342 6476 868 6486
rect 970 6456 1500 6466
rect 970 6390 980 6456
rect 1490 6390 1500 6456
rect 970 6380 1500 6390
rect 342 6360 868 6370
rect 342 6294 352 6360
rect 858 6294 868 6360
rect 342 6284 868 6294
rect 970 6264 1500 6274
rect 970 6198 980 6264
rect 1490 6198 1500 6264
rect 970 6188 1500 6198
rect 342 6168 868 6178
rect 342 6102 352 6168
rect 858 6102 868 6168
rect 342 6092 868 6102
rect 970 6072 1500 6082
rect 970 6006 980 6072
rect 1490 6006 1500 6072
rect 970 5996 1500 6006
rect 342 5976 868 5986
rect 342 5910 352 5976
rect 858 5910 868 5976
rect 342 5900 868 5910
rect 970 5880 1500 5890
rect 970 5814 980 5880
rect 1490 5814 1500 5880
rect 970 5804 1500 5814
rect 342 5784 868 5794
rect 342 5718 352 5784
rect 858 5718 868 5784
rect 342 5708 868 5718
rect 970 5688 1500 5698
rect 970 5622 980 5688
rect 1490 5622 1500 5688
rect 970 5612 1500 5622
rect 342 5592 868 5602
rect 342 5526 352 5592
rect 858 5526 868 5592
rect 342 5516 868 5526
rect 970 5496 1500 5506
rect 970 5430 980 5496
rect 1490 5430 1500 5496
rect 970 5420 1500 5430
rect 342 5400 868 5410
rect 342 5334 352 5400
rect 858 5334 868 5400
rect 342 5324 868 5334
rect 970 5304 1500 5314
rect 970 5238 980 5304
rect 1490 5238 1500 5304
rect 970 5228 1500 5238
rect 342 5208 868 5218
rect 342 5142 352 5208
rect 858 5142 868 5208
rect 342 5132 868 5142
rect 970 5112 1500 5122
rect 970 5046 980 5112
rect 1490 5046 1500 5112
rect 970 5036 1500 5046
rect 342 5016 868 5026
rect 342 4950 352 5016
rect 858 4950 868 5016
rect 342 4940 868 4950
rect 970 4920 1500 4930
rect 970 4854 980 4920
rect 1490 4854 1500 4920
rect 970 4844 1500 4854
rect 342 4824 868 4834
rect 342 4758 352 4824
rect 858 4758 868 4824
rect 342 4748 868 4758
rect 970 4728 1500 4738
rect 970 4662 980 4728
rect 1490 4662 1500 4728
rect 970 4652 1500 4662
rect 342 4632 868 4642
rect 342 4566 352 4632
rect 858 4566 868 4632
rect 342 4556 868 4566
rect 970 4536 1500 4546
rect 970 4470 980 4536
rect 1490 4470 1500 4536
rect 970 4460 1500 4470
rect 342 4440 868 4450
rect 342 4374 352 4440
rect 858 4374 868 4440
rect 342 4364 868 4374
rect 970 4344 1500 4354
rect 970 4278 980 4344
rect 1490 4278 1500 4344
rect 970 4268 1500 4278
rect 342 4248 868 4258
rect 342 4182 352 4248
rect 858 4182 868 4248
rect 342 4172 868 4182
rect 970 4152 1500 4162
rect 970 4086 980 4152
rect 1490 4086 1500 4152
rect 970 4076 1500 4086
rect 342 4056 868 4066
rect 342 3990 352 4056
rect 858 3990 868 4056
rect 342 3980 868 3990
rect 970 3960 1500 3970
rect 970 3894 980 3960
rect 1490 3894 1500 3960
rect 970 3884 1500 3894
rect 342 3864 868 3874
rect 342 3798 352 3864
rect 858 3798 868 3864
rect 342 3788 868 3798
rect 970 3768 1500 3778
rect 970 3702 980 3768
rect 1490 3702 1500 3768
rect 970 3692 1500 3702
rect 342 3672 868 3682
rect 342 3606 352 3672
rect 858 3606 868 3672
rect 342 3596 868 3606
rect 970 3576 1500 3586
rect 970 3510 980 3576
rect 1490 3510 1500 3576
rect 970 3500 1500 3510
rect 342 3480 868 3490
rect 342 3414 352 3480
rect 858 3414 868 3480
rect 342 3404 868 3414
rect 970 3384 1500 3394
rect 970 3318 980 3384
rect 1490 3318 1500 3384
rect 970 3308 1500 3318
rect 342 3288 868 3298
rect 342 3222 352 3288
rect 858 3222 868 3288
rect 342 3212 868 3222
rect 970 3192 1500 3202
rect 970 3126 980 3192
rect 1490 3126 1500 3192
rect 970 3116 1500 3126
rect 342 3096 868 3106
rect 342 3030 352 3096
rect 858 3030 868 3096
rect 342 3020 868 3030
rect 970 3000 1500 3010
rect 970 2934 980 3000
rect 1490 2934 1500 3000
rect 970 2924 1500 2934
rect 342 2904 868 2914
rect 342 2838 352 2904
rect 858 2838 868 2904
rect 342 2828 868 2838
rect 970 2808 1500 2818
rect 970 2742 980 2808
rect 1490 2742 1500 2808
rect 970 2732 1500 2742
rect 342 2712 868 2722
rect 342 2646 352 2712
rect 858 2646 868 2712
rect 342 2636 868 2646
rect 970 2616 1500 2626
rect 970 2550 980 2616
rect 1490 2550 1500 2616
rect 970 2540 1500 2550
rect 342 2520 868 2530
rect 342 2454 352 2520
rect 858 2454 868 2520
rect 342 2444 868 2454
rect 970 2424 1500 2434
rect 970 2358 980 2424
rect 1490 2358 1500 2424
rect 970 2348 1500 2358
rect 342 2328 868 2338
rect 342 2262 352 2328
rect 858 2262 868 2328
rect 342 2252 868 2262
rect 970 2232 1500 2242
rect 970 2166 980 2232
rect 1490 2166 1500 2232
rect 970 2156 1500 2166
rect 342 2136 868 2146
rect 342 2070 352 2136
rect 858 2070 868 2136
rect 342 2060 868 2070
rect 970 2040 1500 2050
rect 970 1974 980 2040
rect 1490 1974 1500 2040
rect 970 1964 1500 1974
rect 342 1944 868 1954
rect 342 1878 352 1944
rect 858 1878 868 1944
rect 342 1868 868 1878
rect 970 1848 1500 1858
rect 970 1782 980 1848
rect 1490 1782 1500 1848
rect 970 1772 1500 1782
rect 342 1752 868 1762
rect 342 1686 352 1752
rect 858 1686 868 1752
rect 342 1676 868 1686
rect 970 1656 1500 1666
rect 970 1590 980 1656
rect 1490 1590 1500 1656
rect 970 1580 1500 1590
rect 342 1560 868 1570
rect 342 1494 352 1560
rect 858 1494 868 1560
rect 342 1484 868 1494
rect 970 1464 1500 1474
rect 970 1398 980 1464
rect 1490 1398 1500 1464
rect 970 1388 1500 1398
rect 342 1368 868 1378
rect 342 1302 352 1368
rect 858 1302 868 1368
rect 342 1292 868 1302
rect 970 1272 1500 1282
rect 970 1206 980 1272
rect 1490 1206 1500 1272
rect 970 1196 1500 1206
rect 342 1176 868 1186
rect 342 1110 352 1176
rect 858 1110 868 1176
rect 342 1100 868 1110
rect 970 1080 1500 1090
rect 970 1014 980 1080
rect 1490 1014 1500 1080
rect 970 1004 1500 1014
rect 342 984 868 994
rect 342 918 352 984
rect 858 918 868 984
rect 342 908 868 918
rect 970 888 1500 898
rect 970 822 980 888
rect 1490 822 1500 888
rect 970 812 1500 822
rect 342 792 868 802
rect 342 726 352 792
rect 858 726 868 792
rect 342 716 868 726
rect 970 696 1500 706
rect 970 630 980 696
rect 1490 630 1500 696
rect 970 620 1500 630
rect 342 600 868 610
rect 342 534 352 600
rect 858 534 868 600
rect 342 524 868 534
<< via3 >>
rect 132 45062 1706 45136
rect 352 44152 858 44218
rect 980 44056 1490 44122
rect 352 43960 858 44026
rect 980 43864 1490 43930
rect 352 43768 858 43834
rect 980 43672 1490 43738
rect 352 43576 858 43642
rect 980 43480 1490 43546
rect 352 43384 858 43450
rect 980 43288 1490 43354
rect 352 43192 858 43258
rect 980 43096 1490 43162
rect 352 43000 858 43066
rect 980 42904 1490 42970
rect 352 42808 858 42874
rect 980 42712 1490 42778
rect 352 42616 858 42682
rect 980 42520 1490 42586
rect 352 42424 858 42490
rect 980 42328 1490 42394
rect 352 42232 858 42298
rect 980 42136 1490 42202
rect 352 42040 858 42106
rect 980 41944 1490 42010
rect 352 41848 858 41914
rect 980 41752 1490 41818
rect 352 41656 858 41722
rect 980 41560 1490 41626
rect 352 41464 858 41530
rect 980 41368 1490 41434
rect 352 41272 858 41338
rect 980 41176 1490 41242
rect 352 41080 858 41146
rect 980 40984 1490 41050
rect 352 40888 858 40954
rect 980 40792 1490 40858
rect 352 40696 858 40762
rect 980 40600 1490 40666
rect 352 40504 858 40570
rect 980 40408 1490 40474
rect 352 40312 858 40378
rect 980 40216 1490 40282
rect 352 40120 858 40186
rect 980 40024 1490 40090
rect 352 39928 858 39994
rect 980 39832 1490 39898
rect 352 39736 858 39802
rect 980 39640 1490 39706
rect 352 39544 858 39610
rect 980 39448 1490 39514
rect 352 39352 858 39418
rect 980 39256 1490 39322
rect 352 39160 858 39226
rect 980 39064 1490 39130
rect 352 38968 858 39034
rect 980 38872 1490 38938
rect 352 38776 858 38842
rect 980 38680 1490 38746
rect 352 38584 858 38650
rect 980 38488 1490 38554
rect 352 38392 858 38458
rect 980 38296 1490 38362
rect 352 38200 858 38266
rect 980 38104 1490 38170
rect 352 38008 858 38074
rect 980 37912 1490 37978
rect 352 37816 858 37882
rect 980 37720 1490 37786
rect 352 37624 858 37690
rect 980 37528 1490 37594
rect 352 37432 858 37498
rect 980 37336 1490 37402
rect 352 37240 858 37306
rect 980 37144 1490 37210
rect 352 37048 858 37114
rect 980 36952 1490 37018
rect 352 36856 858 36922
rect 980 36760 1490 36826
rect 352 36664 858 36730
rect 980 36568 1490 36634
rect 352 36472 858 36538
rect 980 36376 1490 36442
rect 352 36280 858 36346
rect 980 36184 1490 36250
rect 352 36088 858 36154
rect 980 35992 1490 36058
rect 352 35896 858 35962
rect 980 35800 1490 35866
rect 352 35704 858 35770
rect 980 35608 1490 35674
rect 352 35512 858 35578
rect 980 35416 1490 35482
rect 352 35320 858 35386
rect 980 35224 1490 35290
rect 352 35128 858 35194
rect 980 35032 1490 35098
rect 352 34936 858 35002
rect 980 34840 1490 34906
rect 352 34744 858 34810
rect 980 34648 1490 34714
rect 352 34552 858 34618
rect 980 34456 1490 34522
rect 352 34360 858 34426
rect 980 34264 1490 34330
rect 352 34168 858 34234
rect 980 34072 1490 34138
rect 352 33976 858 34042
rect 980 33880 1490 33946
rect 352 33784 858 33850
rect 980 33688 1490 33754
rect 352 33592 858 33658
rect 980 33496 1490 33562
rect 352 33400 858 33466
rect 980 33304 1490 33370
rect 352 33208 858 33274
rect 980 33112 1490 33178
rect 352 33016 858 33082
rect 980 32920 1490 32986
rect 352 32824 858 32890
rect 980 32728 1490 32794
rect 352 32632 858 32698
rect 980 32536 1490 32602
rect 352 32440 858 32506
rect 980 32344 1490 32410
rect 352 32248 858 32314
rect 980 32152 1490 32218
rect 352 32056 858 32122
rect 980 31960 1490 32026
rect 352 31864 858 31930
rect 980 31768 1490 31834
rect 352 31672 858 31738
rect 980 31576 1490 31642
rect 352 31480 858 31546
rect 980 31384 1490 31450
rect 352 31288 858 31354
rect 980 31192 1490 31258
rect 352 31096 858 31162
rect 980 31000 1490 31066
rect 352 30904 858 30970
rect 980 30808 1490 30874
rect 352 30712 858 30778
rect 980 30616 1490 30682
rect 352 30520 858 30586
rect 980 30424 1490 30490
rect 352 30328 858 30394
rect 980 30232 1490 30298
rect 352 30136 858 30202
rect 980 30040 1490 30106
rect 352 29944 858 30010
rect 980 29848 1490 29914
rect 352 29752 858 29818
rect 980 29656 1490 29722
rect 352 29560 858 29626
rect 980 29464 1490 29530
rect 352 29368 858 29434
rect 980 29272 1490 29338
rect 352 29176 858 29242
rect 980 29080 1490 29146
rect 352 28984 858 29050
rect 980 28888 1490 28954
rect 352 28792 858 28858
rect 980 28696 1490 28762
rect 352 28600 858 28666
rect 980 28504 1490 28570
rect 352 28408 858 28474
rect 980 28312 1490 28378
rect 352 28216 858 28282
rect 980 28120 1490 28186
rect 352 28024 858 28090
rect 980 27928 1490 27994
rect 352 27832 858 27898
rect 980 27736 1490 27802
rect 352 27640 858 27706
rect 980 27544 1490 27610
rect 352 27448 858 27514
rect 980 27352 1490 27418
rect 352 27256 858 27322
rect 980 27160 1490 27226
rect 352 27064 858 27130
rect 980 26968 1490 27034
rect 352 26872 858 26938
rect 980 26776 1490 26842
rect 352 26680 858 26746
rect 980 26584 1490 26650
rect 352 26488 858 26554
rect 980 26392 1490 26458
rect 352 26296 858 26362
rect 980 26200 1490 26266
rect 352 26104 858 26170
rect 980 26008 1490 26074
rect 352 25912 858 25978
rect 980 25816 1490 25882
rect 352 25720 858 25786
rect 980 25624 1490 25690
rect 352 25528 858 25594
rect 980 25432 1490 25498
rect 352 25336 858 25402
rect 980 25240 1490 25306
rect 352 25144 858 25210
rect 980 25048 1490 25114
rect 352 24952 858 25018
rect 980 24856 1490 24922
rect 352 24760 858 24826
rect 980 24664 1490 24730
rect 352 24568 858 24634
rect 980 24472 1490 24538
rect 352 24376 858 24442
rect 980 24280 1490 24346
rect 352 24184 858 24250
rect 980 24088 1490 24154
rect 352 23992 858 24058
rect 980 23896 1490 23962
rect 352 23800 858 23866
rect 980 23704 1490 23770
rect 352 23608 858 23674
rect 980 23512 1490 23578
rect 352 23416 858 23482
rect 980 23320 1490 23386
rect 352 23224 858 23290
rect 980 23128 1490 23194
rect 352 23032 858 23098
rect 340 21986 870 22768
rect 352 21654 858 21720
rect 980 21558 1490 21624
rect 352 21462 858 21528
rect 980 21366 1490 21432
rect 352 21270 858 21336
rect 980 21174 1490 21240
rect 352 21078 858 21144
rect 980 20982 1490 21048
rect 352 20886 858 20952
rect 980 20790 1490 20856
rect 352 20694 858 20760
rect 980 20598 1490 20664
rect 352 20502 858 20568
rect 980 20406 1490 20472
rect 352 20310 858 20376
rect 980 20214 1490 20280
rect 352 20118 858 20184
rect 980 20022 1490 20088
rect 352 19926 858 19992
rect 980 19830 1490 19896
rect 352 19734 858 19800
rect 980 19638 1490 19704
rect 352 19542 858 19608
rect 980 19446 1490 19512
rect 352 19350 858 19416
rect 980 19254 1490 19320
rect 352 19158 858 19224
rect 980 19062 1490 19128
rect 352 18966 858 19032
rect 980 18870 1490 18936
rect 352 18774 858 18840
rect 980 18678 1490 18744
rect 352 18582 858 18648
rect 980 18486 1490 18552
rect 352 18390 858 18456
rect 980 18294 1490 18360
rect 352 18198 858 18264
rect 980 18102 1490 18168
rect 352 18006 858 18072
rect 980 17910 1490 17976
rect 352 17814 858 17880
rect 980 17718 1490 17784
rect 352 17622 858 17688
rect 980 17526 1490 17592
rect 352 17430 858 17496
rect 980 17334 1490 17400
rect 352 17238 858 17304
rect 980 17142 1490 17208
rect 352 17046 858 17112
rect 980 16950 1490 17016
rect 352 16854 858 16920
rect 980 16758 1490 16824
rect 352 16662 858 16728
rect 980 16566 1490 16632
rect 352 16470 858 16536
rect 980 16374 1490 16440
rect 352 16278 858 16344
rect 980 16182 1490 16248
rect 352 16086 858 16152
rect 980 15990 1490 16056
rect 352 15894 858 15960
rect 980 15798 1490 15864
rect 352 15702 858 15768
rect 980 15606 1490 15672
rect 352 15510 858 15576
rect 980 15414 1490 15480
rect 352 15318 858 15384
rect 980 15222 1490 15288
rect 352 15126 858 15192
rect 980 15030 1490 15096
rect 352 14934 858 15000
rect 980 14838 1490 14904
rect 352 14742 858 14808
rect 980 14646 1490 14712
rect 352 14550 858 14616
rect 980 14454 1490 14520
rect 352 14358 858 14424
rect 980 14262 1490 14328
rect 352 14166 858 14232
rect 980 14070 1490 14136
rect 352 13974 858 14040
rect 980 13878 1490 13944
rect 352 13782 858 13848
rect 980 13686 1490 13752
rect 352 13590 858 13656
rect 980 13494 1490 13560
rect 352 13398 858 13464
rect 980 13302 1490 13368
rect 352 13206 858 13272
rect 980 13110 1490 13176
rect 352 13014 858 13080
rect 980 12918 1490 12984
rect 352 12822 858 12888
rect 980 12726 1490 12792
rect 352 12630 858 12696
rect 980 12534 1490 12600
rect 352 12438 858 12504
rect 980 12342 1490 12408
rect 352 12246 858 12312
rect 980 12150 1490 12216
rect 352 12054 858 12120
rect 980 11958 1490 12024
rect 352 11862 858 11928
rect 980 11766 1490 11832
rect 352 11670 858 11736
rect 980 11574 1490 11640
rect 352 11478 858 11544
rect 980 11382 1490 11448
rect 352 11286 858 11352
rect 980 11190 1490 11256
rect 352 11094 858 11160
rect 980 10998 1490 11064
rect 352 10902 858 10968
rect 980 10806 1490 10872
rect 352 10710 858 10776
rect 980 10614 1490 10680
rect 352 10518 858 10584
rect 980 10422 1490 10488
rect 352 10326 858 10392
rect 980 10230 1490 10296
rect 352 10134 858 10200
rect 980 10038 1490 10104
rect 352 9942 858 10008
rect 980 9846 1490 9912
rect 352 9750 858 9816
rect 980 9654 1490 9720
rect 352 9558 858 9624
rect 980 9462 1490 9528
rect 352 9366 858 9432
rect 980 9270 1490 9336
rect 352 9174 858 9240
rect 980 9078 1490 9144
rect 352 8982 858 9048
rect 980 8886 1490 8952
rect 352 8790 858 8856
rect 980 8694 1490 8760
rect 352 8598 858 8664
rect 980 8502 1490 8568
rect 352 8406 858 8472
rect 980 8310 1490 8376
rect 352 8214 858 8280
rect 980 8118 1490 8184
rect 352 8022 858 8088
rect 980 7926 1490 7992
rect 352 7830 858 7896
rect 980 7734 1490 7800
rect 352 7638 858 7704
rect 980 7542 1490 7608
rect 352 7446 858 7512
rect 980 7350 1490 7416
rect 352 7254 858 7320
rect 980 7158 1490 7224
rect 352 7062 858 7128
rect 980 6966 1490 7032
rect 352 6870 858 6936
rect 980 6774 1490 6840
rect 352 6678 858 6744
rect 980 6582 1490 6648
rect 352 6486 858 6552
rect 980 6390 1490 6456
rect 352 6294 858 6360
rect 980 6198 1490 6264
rect 352 6102 858 6168
rect 980 6006 1490 6072
rect 352 5910 858 5976
rect 980 5814 1490 5880
rect 352 5718 858 5784
rect 980 5622 1490 5688
rect 352 5526 858 5592
rect 980 5430 1490 5496
rect 352 5334 858 5400
rect 980 5238 1490 5304
rect 352 5142 858 5208
rect 980 5046 1490 5112
rect 352 4950 858 5016
rect 980 4854 1490 4920
rect 352 4758 858 4824
rect 980 4662 1490 4728
rect 352 4566 858 4632
rect 980 4470 1490 4536
rect 352 4374 858 4440
rect 980 4278 1490 4344
rect 352 4182 858 4248
rect 980 4086 1490 4152
rect 352 3990 858 4056
rect 980 3894 1490 3960
rect 352 3798 858 3864
rect 980 3702 1490 3768
rect 352 3606 858 3672
rect 980 3510 1490 3576
rect 352 3414 858 3480
rect 980 3318 1490 3384
rect 352 3222 858 3288
rect 980 3126 1490 3192
rect 352 3030 858 3096
rect 980 2934 1490 3000
rect 352 2838 858 2904
rect 980 2742 1490 2808
rect 352 2646 858 2712
rect 980 2550 1490 2616
rect 352 2454 858 2520
rect 980 2358 1490 2424
rect 352 2262 858 2328
rect 980 2166 1490 2232
rect 352 2070 858 2136
rect 980 1974 1490 2040
rect 352 1878 858 1944
rect 980 1782 1490 1848
rect 352 1686 858 1752
rect 980 1590 1490 1656
rect 352 1494 858 1560
rect 980 1398 1490 1464
rect 352 1302 858 1368
rect 980 1206 1490 1272
rect 352 1110 858 1176
rect 980 1014 1490 1080
rect 352 918 858 984
rect 980 822 1490 888
rect 352 726 858 792
rect 980 630 1490 696
rect 352 534 858 600
<< metal4 >>
rect 0 45136 1840 45152
rect 0 45062 132 45136
rect 1706 45062 1840 45136
rect 0 45052 1840 45062
rect 0 0 240 44848
rect 340 44218 870 44848
rect 340 44152 352 44218
rect 858 44152 870 44218
rect 340 44026 870 44152
rect 340 43960 352 44026
rect 858 43960 870 44026
rect 340 43834 870 43960
rect 340 43768 352 43834
rect 858 43768 870 43834
rect 340 43642 870 43768
rect 340 43576 352 43642
rect 858 43576 870 43642
rect 340 43450 870 43576
rect 340 43384 352 43450
rect 858 43384 870 43450
rect 340 43258 870 43384
rect 340 43192 352 43258
rect 858 43192 870 43258
rect 340 43066 870 43192
rect 340 43000 352 43066
rect 858 43000 870 43066
rect 340 42874 870 43000
rect 340 42808 352 42874
rect 858 42808 870 42874
rect 340 42682 870 42808
rect 340 42616 352 42682
rect 858 42616 870 42682
rect 340 42490 870 42616
rect 340 42424 352 42490
rect 858 42424 870 42490
rect 340 42298 870 42424
rect 340 42232 352 42298
rect 858 42232 870 42298
rect 340 42106 870 42232
rect 340 42040 352 42106
rect 858 42040 870 42106
rect 340 41914 870 42040
rect 340 41848 352 41914
rect 858 41848 870 41914
rect 340 41722 870 41848
rect 340 41656 352 41722
rect 858 41656 870 41722
rect 340 41530 870 41656
rect 340 41464 352 41530
rect 858 41464 870 41530
rect 340 41338 870 41464
rect 340 41272 352 41338
rect 858 41272 870 41338
rect 340 41146 870 41272
rect 340 41080 352 41146
rect 858 41080 870 41146
rect 340 40954 870 41080
rect 340 40888 352 40954
rect 858 40888 870 40954
rect 340 40762 870 40888
rect 340 40696 352 40762
rect 858 40696 870 40762
rect 340 40570 870 40696
rect 340 40504 352 40570
rect 858 40504 870 40570
rect 340 40378 870 40504
rect 340 40312 352 40378
rect 858 40312 870 40378
rect 340 40186 870 40312
rect 340 40120 352 40186
rect 858 40120 870 40186
rect 340 39994 870 40120
rect 340 39928 352 39994
rect 858 39928 870 39994
rect 340 39802 870 39928
rect 340 39736 352 39802
rect 858 39736 870 39802
rect 340 39610 870 39736
rect 340 39544 352 39610
rect 858 39544 870 39610
rect 340 39418 870 39544
rect 340 39352 352 39418
rect 858 39352 870 39418
rect 340 39226 870 39352
rect 340 39160 352 39226
rect 858 39160 870 39226
rect 340 39034 870 39160
rect 340 38968 352 39034
rect 858 38968 870 39034
rect 340 38842 870 38968
rect 340 38776 352 38842
rect 858 38776 870 38842
rect 340 38650 870 38776
rect 340 38584 352 38650
rect 858 38584 870 38650
rect 340 38458 870 38584
rect 340 38392 352 38458
rect 858 38392 870 38458
rect 340 38266 870 38392
rect 340 38200 352 38266
rect 858 38200 870 38266
rect 340 38074 870 38200
rect 340 38008 352 38074
rect 858 38008 870 38074
rect 340 37882 870 38008
rect 340 37816 352 37882
rect 858 37816 870 37882
rect 340 37690 870 37816
rect 340 37624 352 37690
rect 858 37624 870 37690
rect 340 37498 870 37624
rect 340 37432 352 37498
rect 858 37432 870 37498
rect 340 37306 870 37432
rect 340 37240 352 37306
rect 858 37240 870 37306
rect 340 37114 870 37240
rect 340 37048 352 37114
rect 858 37048 870 37114
rect 340 36922 870 37048
rect 340 36856 352 36922
rect 858 36856 870 36922
rect 340 36730 870 36856
rect 340 36664 352 36730
rect 858 36664 870 36730
rect 340 36538 870 36664
rect 340 36472 352 36538
rect 858 36472 870 36538
rect 340 36346 870 36472
rect 340 36280 352 36346
rect 858 36280 870 36346
rect 340 36154 870 36280
rect 340 36088 352 36154
rect 858 36088 870 36154
rect 340 35962 870 36088
rect 340 35896 352 35962
rect 858 35896 870 35962
rect 340 35770 870 35896
rect 340 35704 352 35770
rect 858 35704 870 35770
rect 340 35578 870 35704
rect 340 35512 352 35578
rect 858 35512 870 35578
rect 340 35386 870 35512
rect 340 35320 352 35386
rect 858 35320 870 35386
rect 340 35194 870 35320
rect 340 35128 352 35194
rect 858 35128 870 35194
rect 340 35002 870 35128
rect 340 34936 352 35002
rect 858 34936 870 35002
rect 340 34810 870 34936
rect 340 34744 352 34810
rect 858 34744 870 34810
rect 340 34618 870 34744
rect 340 34552 352 34618
rect 858 34552 870 34618
rect 340 34426 870 34552
rect 340 34360 352 34426
rect 858 34360 870 34426
rect 340 34234 870 34360
rect 340 34168 352 34234
rect 858 34168 870 34234
rect 340 34042 870 34168
rect 340 33976 352 34042
rect 858 33976 870 34042
rect 340 33850 870 33976
rect 340 33784 352 33850
rect 858 33784 870 33850
rect 340 33658 870 33784
rect 340 33592 352 33658
rect 858 33592 870 33658
rect 340 33466 870 33592
rect 340 33400 352 33466
rect 858 33400 870 33466
rect 340 33274 870 33400
rect 340 33208 352 33274
rect 858 33208 870 33274
rect 340 33082 870 33208
rect 340 33016 352 33082
rect 858 33016 870 33082
rect 340 32890 870 33016
rect 340 32824 352 32890
rect 858 32824 870 32890
rect 340 32698 870 32824
rect 340 32632 352 32698
rect 858 32632 870 32698
rect 340 32506 870 32632
rect 340 32440 352 32506
rect 858 32440 870 32506
rect 340 32314 870 32440
rect 340 32248 352 32314
rect 858 32248 870 32314
rect 340 32122 870 32248
rect 340 32056 352 32122
rect 858 32056 870 32122
rect 340 31930 870 32056
rect 340 31864 352 31930
rect 858 31864 870 31930
rect 340 31738 870 31864
rect 340 31672 352 31738
rect 858 31672 870 31738
rect 340 31546 870 31672
rect 340 31480 352 31546
rect 858 31480 870 31546
rect 340 31354 870 31480
rect 340 31288 352 31354
rect 858 31288 870 31354
rect 340 31162 870 31288
rect 340 31096 352 31162
rect 858 31096 870 31162
rect 340 30970 870 31096
rect 340 30904 352 30970
rect 858 30904 870 30970
rect 340 30778 870 30904
rect 340 30712 352 30778
rect 858 30712 870 30778
rect 340 30586 870 30712
rect 340 30520 352 30586
rect 858 30520 870 30586
rect 340 30394 870 30520
rect 340 30328 352 30394
rect 858 30328 870 30394
rect 340 30202 870 30328
rect 340 30136 352 30202
rect 858 30136 870 30202
rect 340 30010 870 30136
rect 340 29944 352 30010
rect 858 29944 870 30010
rect 340 29818 870 29944
rect 340 29752 352 29818
rect 858 29752 870 29818
rect 340 29626 870 29752
rect 340 29560 352 29626
rect 858 29560 870 29626
rect 340 29434 870 29560
rect 340 29368 352 29434
rect 858 29368 870 29434
rect 340 29242 870 29368
rect 340 29176 352 29242
rect 858 29176 870 29242
rect 340 29050 870 29176
rect 340 28984 352 29050
rect 858 28984 870 29050
rect 340 28858 870 28984
rect 340 28792 352 28858
rect 858 28792 870 28858
rect 340 28666 870 28792
rect 340 28600 352 28666
rect 858 28600 870 28666
rect 340 28474 870 28600
rect 340 28408 352 28474
rect 858 28408 870 28474
rect 340 28282 870 28408
rect 340 28216 352 28282
rect 858 28216 870 28282
rect 340 28090 870 28216
rect 340 28024 352 28090
rect 858 28024 870 28090
rect 340 27898 870 28024
rect 340 27832 352 27898
rect 858 27832 870 27898
rect 340 27706 870 27832
rect 340 27640 352 27706
rect 858 27640 870 27706
rect 340 27514 870 27640
rect 340 27448 352 27514
rect 858 27448 870 27514
rect 340 27322 870 27448
rect 340 27256 352 27322
rect 858 27256 870 27322
rect 340 27130 870 27256
rect 340 27064 352 27130
rect 858 27064 870 27130
rect 340 26938 870 27064
rect 340 26872 352 26938
rect 858 26872 870 26938
rect 340 26746 870 26872
rect 340 26680 352 26746
rect 858 26680 870 26746
rect 340 26554 870 26680
rect 340 26488 352 26554
rect 858 26488 870 26554
rect 340 26362 870 26488
rect 340 26296 352 26362
rect 858 26296 870 26362
rect 340 26170 870 26296
rect 340 26104 352 26170
rect 858 26104 870 26170
rect 340 25978 870 26104
rect 340 25912 352 25978
rect 858 25912 870 25978
rect 340 25786 870 25912
rect 340 25720 352 25786
rect 858 25720 870 25786
rect 340 25594 870 25720
rect 340 25528 352 25594
rect 858 25528 870 25594
rect 340 25402 870 25528
rect 340 25336 352 25402
rect 858 25336 870 25402
rect 340 25210 870 25336
rect 340 25144 352 25210
rect 858 25144 870 25210
rect 340 25018 870 25144
rect 340 24952 352 25018
rect 858 24952 870 25018
rect 340 24826 870 24952
rect 340 24760 352 24826
rect 858 24760 870 24826
rect 340 24634 870 24760
rect 340 24568 352 24634
rect 858 24568 870 24634
rect 340 24497 870 24568
rect 970 44122 1500 44848
rect 970 44056 980 44122
rect 1490 44056 1500 44122
rect 970 43930 1500 44056
rect 970 43864 980 43930
rect 1490 43864 1500 43930
rect 970 43738 1500 43864
rect 970 43672 980 43738
rect 1490 43672 1500 43738
rect 970 43546 1500 43672
rect 970 43480 980 43546
rect 1490 43480 1500 43546
rect 970 43354 1500 43480
rect 970 43288 980 43354
rect 1490 43288 1500 43354
rect 970 43162 1500 43288
rect 970 43096 980 43162
rect 1490 43096 1500 43162
rect 970 42970 1500 43096
rect 970 42904 980 42970
rect 1490 42904 1500 42970
rect 970 42778 1500 42904
rect 970 42712 980 42778
rect 1490 42712 1500 42778
rect 970 42586 1500 42712
rect 970 42520 980 42586
rect 1490 42520 1500 42586
rect 970 42394 1500 42520
rect 970 42328 980 42394
rect 1490 42328 1500 42394
rect 970 42202 1500 42328
rect 970 42136 980 42202
rect 1490 42136 1500 42202
rect 970 42010 1500 42136
rect 970 41944 980 42010
rect 1490 41944 1500 42010
rect 970 41818 1500 41944
rect 970 41752 980 41818
rect 1490 41752 1500 41818
rect 970 41626 1500 41752
rect 970 41560 980 41626
rect 1490 41560 1500 41626
rect 970 41434 1500 41560
rect 970 41368 980 41434
rect 1490 41368 1500 41434
rect 970 41242 1500 41368
rect 970 41176 980 41242
rect 1490 41176 1500 41242
rect 970 41050 1500 41176
rect 970 40984 980 41050
rect 1490 40984 1500 41050
rect 970 40858 1500 40984
rect 970 40792 980 40858
rect 1490 40792 1500 40858
rect 970 40666 1500 40792
rect 970 40600 980 40666
rect 1490 40600 1500 40666
rect 970 40474 1500 40600
rect 970 40408 980 40474
rect 1490 40408 1500 40474
rect 970 40282 1500 40408
rect 970 40216 980 40282
rect 1490 40216 1500 40282
rect 970 40090 1500 40216
rect 970 40024 980 40090
rect 1490 40024 1500 40090
rect 970 39898 1500 40024
rect 970 39832 980 39898
rect 1490 39832 1500 39898
rect 970 39706 1500 39832
rect 970 39640 980 39706
rect 1490 39640 1500 39706
rect 970 39514 1500 39640
rect 970 39448 980 39514
rect 1490 39448 1500 39514
rect 970 39322 1500 39448
rect 970 39256 980 39322
rect 1490 39256 1500 39322
rect 970 39130 1500 39256
rect 970 39064 980 39130
rect 1490 39064 1500 39130
rect 970 38938 1500 39064
rect 970 38872 980 38938
rect 1490 38872 1500 38938
rect 970 38746 1500 38872
rect 970 38680 980 38746
rect 1490 38680 1500 38746
rect 970 38554 1500 38680
rect 970 38488 980 38554
rect 1490 38488 1500 38554
rect 970 38362 1500 38488
rect 970 38296 980 38362
rect 1490 38296 1500 38362
rect 970 38170 1500 38296
rect 970 38104 980 38170
rect 1490 38104 1500 38170
rect 970 37978 1500 38104
rect 970 37912 980 37978
rect 1490 37912 1500 37978
rect 970 37786 1500 37912
rect 970 37720 980 37786
rect 1490 37720 1500 37786
rect 970 37594 1500 37720
rect 970 37528 980 37594
rect 1490 37528 1500 37594
rect 970 37402 1500 37528
rect 970 37336 980 37402
rect 1490 37336 1500 37402
rect 970 37210 1500 37336
rect 970 37144 980 37210
rect 1490 37144 1500 37210
rect 970 37018 1500 37144
rect 970 36952 980 37018
rect 1490 36952 1500 37018
rect 970 36826 1500 36952
rect 970 36760 980 36826
rect 1490 36760 1500 36826
rect 970 36634 1500 36760
rect 970 36568 980 36634
rect 1490 36568 1500 36634
rect 970 36442 1500 36568
rect 970 36376 980 36442
rect 1490 36376 1500 36442
rect 970 36250 1500 36376
rect 970 36184 980 36250
rect 1490 36184 1500 36250
rect 970 36058 1500 36184
rect 970 35992 980 36058
rect 1490 35992 1500 36058
rect 970 35866 1500 35992
rect 970 35800 980 35866
rect 1490 35800 1500 35866
rect 970 35674 1500 35800
rect 970 35608 980 35674
rect 1490 35608 1500 35674
rect 970 35482 1500 35608
rect 970 35416 980 35482
rect 1490 35416 1500 35482
rect 970 35290 1500 35416
rect 970 35224 980 35290
rect 1490 35224 1500 35290
rect 970 35098 1500 35224
rect 970 35032 980 35098
rect 1490 35032 1500 35098
rect 970 34906 1500 35032
rect 970 34840 980 34906
rect 1490 34840 1500 34906
rect 970 34714 1500 34840
rect 970 34648 980 34714
rect 1490 34648 1500 34714
rect 970 34522 1500 34648
rect 970 34456 980 34522
rect 1490 34456 1500 34522
rect 970 34330 1500 34456
rect 970 34264 980 34330
rect 1490 34264 1500 34330
rect 970 34138 1500 34264
rect 970 34072 980 34138
rect 1490 34072 1500 34138
rect 970 33946 1500 34072
rect 970 33880 980 33946
rect 1490 33880 1500 33946
rect 970 33754 1500 33880
rect 970 33688 980 33754
rect 1490 33688 1500 33754
rect 970 33562 1500 33688
rect 970 33496 980 33562
rect 1490 33496 1500 33562
rect 970 33370 1500 33496
rect 970 33304 980 33370
rect 1490 33304 1500 33370
rect 970 33178 1500 33304
rect 970 33112 980 33178
rect 1490 33112 1500 33178
rect 970 32986 1500 33112
rect 970 32920 980 32986
rect 1490 32920 1500 32986
rect 970 32794 1500 32920
rect 970 32728 980 32794
rect 1490 32728 1500 32794
rect 970 32602 1500 32728
rect 970 32536 980 32602
rect 1490 32536 1500 32602
rect 970 32410 1500 32536
rect 970 32344 980 32410
rect 1490 32344 1500 32410
rect 970 32218 1500 32344
rect 970 32152 980 32218
rect 1490 32152 1500 32218
rect 970 32026 1500 32152
rect 970 31960 980 32026
rect 1490 31960 1500 32026
rect 970 31834 1500 31960
rect 970 31768 980 31834
rect 1490 31768 1500 31834
rect 970 31642 1500 31768
rect 970 31576 980 31642
rect 1490 31576 1500 31642
rect 970 31450 1500 31576
rect 970 31384 980 31450
rect 1490 31384 1500 31450
rect 970 31258 1500 31384
rect 970 31192 980 31258
rect 1490 31192 1500 31258
rect 970 31066 1500 31192
rect 970 31000 980 31066
rect 1490 31000 1500 31066
rect 970 30874 1500 31000
rect 970 30808 980 30874
rect 1490 30808 1500 30874
rect 970 30682 1500 30808
rect 970 30616 980 30682
rect 1490 30616 1500 30682
rect 970 30490 1500 30616
rect 970 30424 980 30490
rect 1490 30424 1500 30490
rect 970 30298 1500 30424
rect 970 30232 980 30298
rect 1490 30232 1500 30298
rect 970 30106 1500 30232
rect 970 30040 980 30106
rect 1490 30040 1500 30106
rect 970 29914 1500 30040
rect 970 29848 980 29914
rect 1490 29848 1500 29914
rect 970 29722 1500 29848
rect 970 29656 980 29722
rect 1490 29656 1500 29722
rect 970 29530 1500 29656
rect 970 29464 980 29530
rect 1490 29464 1500 29530
rect 970 29338 1500 29464
rect 970 29272 980 29338
rect 1490 29272 1500 29338
rect 970 29146 1500 29272
rect 970 29080 980 29146
rect 1490 29080 1500 29146
rect 970 28954 1500 29080
rect 970 28888 980 28954
rect 1490 28888 1500 28954
rect 970 28762 1500 28888
rect 970 28696 980 28762
rect 1490 28696 1500 28762
rect 970 28570 1500 28696
rect 970 28504 980 28570
rect 1490 28504 1500 28570
rect 970 28378 1500 28504
rect 970 28312 980 28378
rect 1490 28312 1500 28378
rect 970 28186 1500 28312
rect 970 28120 980 28186
rect 1490 28120 1500 28186
rect 970 27994 1500 28120
rect 970 27928 980 27994
rect 1490 27928 1500 27994
rect 970 27802 1500 27928
rect 970 27736 980 27802
rect 1490 27736 1500 27802
rect 970 27610 1500 27736
rect 970 27544 980 27610
rect 1490 27544 1500 27610
rect 970 27418 1500 27544
rect 970 27352 980 27418
rect 1490 27352 1500 27418
rect 970 27226 1500 27352
rect 970 27160 980 27226
rect 1490 27160 1500 27226
rect 970 27034 1500 27160
rect 970 26968 980 27034
rect 1490 26968 1500 27034
rect 970 26842 1500 26968
rect 970 26776 980 26842
rect 1490 26776 1500 26842
rect 970 26650 1500 26776
rect 970 26584 980 26650
rect 1490 26584 1500 26650
rect 970 26458 1500 26584
rect 970 26392 980 26458
rect 1490 26392 1500 26458
rect 970 26266 1500 26392
rect 970 26200 980 26266
rect 1490 26200 1500 26266
rect 970 26074 1500 26200
rect 970 26008 980 26074
rect 1490 26008 1500 26074
rect 970 25882 1500 26008
rect 970 25816 980 25882
rect 1490 25816 1500 25882
rect 970 25690 1500 25816
rect 970 25624 980 25690
rect 1490 25624 1500 25690
rect 970 25498 1500 25624
rect 970 25432 980 25498
rect 1490 25432 1500 25498
rect 970 25306 1500 25432
rect 970 25240 980 25306
rect 1490 25240 1500 25306
rect 970 25114 1500 25240
rect 970 25048 980 25114
rect 1490 25048 1500 25114
rect 970 24922 1500 25048
rect 970 24856 980 24922
rect 1490 24856 1500 24922
rect 970 24730 1500 24856
rect 970 24664 980 24730
rect 1490 24664 1500 24730
rect 970 24538 1500 24664
rect 339 24442 871 24497
rect 339 24431 352 24442
rect 340 24376 352 24431
rect 858 24431 871 24442
rect 970 24472 980 24538
rect 1490 24472 1500 24538
rect 858 24376 870 24431
rect 340 24307 870 24376
rect 970 24346 1500 24472
rect 339 24250 871 24307
rect 339 24241 352 24250
rect 340 24184 352 24241
rect 858 24241 871 24250
rect 970 24280 980 24346
rect 1490 24280 1500 24346
rect 858 24184 870 24241
rect 340 24113 870 24184
rect 970 24154 1500 24280
rect 339 24058 871 24113
rect 339 24047 352 24058
rect 340 23992 352 24047
rect 858 24047 871 24058
rect 970 24088 980 24154
rect 1490 24088 1500 24154
rect 858 23992 870 24047
rect 340 23923 870 23992
rect 970 23962 1500 24088
rect 339 23866 871 23923
rect 339 23857 352 23866
rect 340 23800 352 23857
rect 858 23857 871 23866
rect 970 23896 980 23962
rect 1490 23896 1500 23962
rect 858 23800 870 23857
rect 340 23731 870 23800
rect 970 23770 1500 23896
rect 339 23674 871 23731
rect 339 23665 352 23674
rect 340 23608 352 23665
rect 858 23665 871 23674
rect 970 23704 980 23770
rect 1490 23704 1500 23770
rect 858 23608 870 23665
rect 340 23537 870 23608
rect 970 23578 1500 23704
rect 339 23482 871 23537
rect 339 23471 352 23482
rect 340 23416 352 23471
rect 858 23471 871 23482
rect 970 23512 980 23578
rect 1490 23512 1500 23578
rect 858 23416 870 23471
rect 340 23347 870 23416
rect 970 23386 1500 23512
rect 339 23290 871 23347
rect 339 23281 352 23290
rect 340 23224 352 23281
rect 858 23281 871 23290
rect 970 23320 980 23386
rect 1490 23320 1500 23386
rect 858 23224 870 23281
rect 340 23155 870 23224
rect 970 23194 1500 23320
rect 339 23098 871 23155
rect 339 23089 352 23098
rect 340 23032 352 23089
rect 858 23089 871 23098
rect 970 23128 980 23194
rect 1490 23128 1500 23194
rect 858 23032 870 23089
rect 340 22769 870 23032
rect 339 22768 871 22769
rect 339 21986 340 22768
rect 870 21986 871 22768
rect 339 21985 871 21986
rect 340 21720 870 21985
rect 340 21654 352 21720
rect 858 21654 870 21720
rect 340 21528 870 21654
rect 340 21462 352 21528
rect 858 21462 870 21528
rect 340 21336 870 21462
rect 340 21270 352 21336
rect 858 21270 870 21336
rect 340 21144 870 21270
rect 340 21078 352 21144
rect 858 21078 870 21144
rect 340 20952 870 21078
rect 340 20886 352 20952
rect 858 20886 870 20952
rect 340 20760 870 20886
rect 340 20694 352 20760
rect 858 20694 870 20760
rect 340 20568 870 20694
rect 340 20502 352 20568
rect 858 20502 870 20568
rect 340 20376 870 20502
rect 340 20310 352 20376
rect 858 20310 870 20376
rect 340 20184 870 20310
rect 340 20118 352 20184
rect 858 20118 870 20184
rect 340 19992 870 20118
rect 340 19926 352 19992
rect 858 19926 870 19992
rect 340 19800 870 19926
rect 340 19734 352 19800
rect 858 19734 870 19800
rect 340 19608 870 19734
rect 340 19542 352 19608
rect 858 19542 870 19608
rect 340 19416 870 19542
rect 340 19350 352 19416
rect 858 19350 870 19416
rect 340 19224 870 19350
rect 340 19158 352 19224
rect 858 19158 870 19224
rect 340 19032 870 19158
rect 340 18966 352 19032
rect 858 18966 870 19032
rect 340 18840 870 18966
rect 340 18774 352 18840
rect 858 18774 870 18840
rect 340 18648 870 18774
rect 340 18582 352 18648
rect 858 18582 870 18648
rect 340 18456 870 18582
rect 340 18390 352 18456
rect 858 18390 870 18456
rect 340 18264 870 18390
rect 340 18198 352 18264
rect 858 18198 870 18264
rect 340 18072 870 18198
rect 340 18006 352 18072
rect 858 18006 870 18072
rect 340 17880 870 18006
rect 340 17814 352 17880
rect 858 17814 870 17880
rect 340 17688 870 17814
rect 340 17622 352 17688
rect 858 17622 870 17688
rect 340 17496 870 17622
rect 340 17430 352 17496
rect 858 17430 870 17496
rect 340 17304 870 17430
rect 340 17238 352 17304
rect 858 17238 870 17304
rect 340 17112 870 17238
rect 340 17046 352 17112
rect 858 17046 870 17112
rect 340 16920 870 17046
rect 340 16854 352 16920
rect 858 16854 870 16920
rect 340 16728 870 16854
rect 340 16662 352 16728
rect 858 16662 870 16728
rect 340 16536 870 16662
rect 340 16470 352 16536
rect 858 16470 870 16536
rect 340 16344 870 16470
rect 340 16278 352 16344
rect 858 16278 870 16344
rect 340 16152 870 16278
rect 340 16086 352 16152
rect 858 16086 870 16152
rect 340 15960 870 16086
rect 340 15894 352 15960
rect 858 15894 870 15960
rect 340 15768 870 15894
rect 340 15702 352 15768
rect 858 15702 870 15768
rect 340 15576 870 15702
rect 340 15510 352 15576
rect 858 15510 870 15576
rect 340 15384 870 15510
rect 340 15318 352 15384
rect 858 15318 870 15384
rect 340 15192 870 15318
rect 340 15126 352 15192
rect 858 15126 870 15192
rect 340 15000 870 15126
rect 340 14934 352 15000
rect 858 14934 870 15000
rect 340 14808 870 14934
rect 340 14742 352 14808
rect 858 14742 870 14808
rect 340 14616 870 14742
rect 340 14550 352 14616
rect 858 14550 870 14616
rect 340 14424 870 14550
rect 340 14358 352 14424
rect 858 14358 870 14424
rect 340 14232 870 14358
rect 340 14166 352 14232
rect 858 14166 870 14232
rect 340 14040 870 14166
rect 340 13974 352 14040
rect 858 13974 870 14040
rect 340 13848 870 13974
rect 340 13782 352 13848
rect 858 13782 870 13848
rect 340 13656 870 13782
rect 340 13590 352 13656
rect 858 13590 870 13656
rect 340 13464 870 13590
rect 340 13398 352 13464
rect 858 13398 870 13464
rect 340 13272 870 13398
rect 340 13206 352 13272
rect 858 13206 870 13272
rect 340 13080 870 13206
rect 340 13014 352 13080
rect 858 13014 870 13080
rect 340 12888 870 13014
rect 340 12822 352 12888
rect 858 12822 870 12888
rect 340 12696 870 12822
rect 340 12630 352 12696
rect 858 12630 870 12696
rect 340 12504 870 12630
rect 340 12438 352 12504
rect 858 12438 870 12504
rect 340 12312 870 12438
rect 340 12246 352 12312
rect 858 12246 870 12312
rect 340 12120 870 12246
rect 340 12054 352 12120
rect 858 12054 870 12120
rect 340 11928 870 12054
rect 340 11862 352 11928
rect 858 11862 870 11928
rect 340 11736 870 11862
rect 340 11670 352 11736
rect 858 11670 870 11736
rect 340 11544 870 11670
rect 340 11478 352 11544
rect 858 11478 870 11544
rect 340 11352 870 11478
rect 340 11286 352 11352
rect 858 11286 870 11352
rect 340 11160 870 11286
rect 340 11094 352 11160
rect 858 11094 870 11160
rect 340 10968 870 11094
rect 340 10902 352 10968
rect 858 10902 870 10968
rect 340 10776 870 10902
rect 340 10710 352 10776
rect 858 10710 870 10776
rect 340 10584 870 10710
rect 340 10518 352 10584
rect 858 10518 870 10584
rect 340 10392 870 10518
rect 340 10326 352 10392
rect 858 10326 870 10392
rect 340 10200 870 10326
rect 340 10134 352 10200
rect 858 10134 870 10200
rect 340 10008 870 10134
rect 340 9942 352 10008
rect 858 9942 870 10008
rect 340 9816 870 9942
rect 340 9750 352 9816
rect 858 9750 870 9816
rect 340 9624 870 9750
rect 340 9558 352 9624
rect 858 9558 870 9624
rect 340 9432 870 9558
rect 340 9366 352 9432
rect 858 9366 870 9432
rect 340 9240 870 9366
rect 340 9174 352 9240
rect 858 9174 870 9240
rect 340 9048 870 9174
rect 340 8982 352 9048
rect 858 8982 870 9048
rect 340 8856 870 8982
rect 340 8790 352 8856
rect 858 8790 870 8856
rect 340 8664 870 8790
rect 340 8598 352 8664
rect 858 8598 870 8664
rect 340 8472 870 8598
rect 340 8406 352 8472
rect 858 8406 870 8472
rect 340 8280 870 8406
rect 340 8214 352 8280
rect 858 8214 870 8280
rect 340 8088 870 8214
rect 340 8022 352 8088
rect 858 8022 870 8088
rect 340 7896 870 8022
rect 340 7830 352 7896
rect 858 7830 870 7896
rect 340 7704 870 7830
rect 340 7638 352 7704
rect 858 7638 870 7704
rect 340 7512 870 7638
rect 340 7446 352 7512
rect 858 7446 870 7512
rect 340 7320 870 7446
rect 340 7254 352 7320
rect 858 7254 870 7320
rect 340 7128 870 7254
rect 340 7062 352 7128
rect 858 7062 870 7128
rect 340 6936 870 7062
rect 340 6870 352 6936
rect 858 6870 870 6936
rect 340 6744 870 6870
rect 340 6678 352 6744
rect 858 6678 870 6744
rect 340 6552 870 6678
rect 340 6486 352 6552
rect 858 6486 870 6552
rect 340 6360 870 6486
rect 340 6294 352 6360
rect 858 6294 870 6360
rect 340 6168 870 6294
rect 340 6102 352 6168
rect 858 6102 870 6168
rect 340 5976 870 6102
rect 340 5910 352 5976
rect 858 5910 870 5976
rect 340 5784 870 5910
rect 340 5718 352 5784
rect 858 5718 870 5784
rect 340 5592 870 5718
rect 340 5526 352 5592
rect 858 5526 870 5592
rect 340 5400 870 5526
rect 340 5334 352 5400
rect 858 5334 870 5400
rect 340 5208 870 5334
rect 340 5142 352 5208
rect 858 5142 870 5208
rect 340 5016 870 5142
rect 340 4950 352 5016
rect 858 4950 870 5016
rect 340 4824 870 4950
rect 340 4758 352 4824
rect 858 4758 870 4824
rect 340 4632 870 4758
rect 340 4566 352 4632
rect 858 4566 870 4632
rect 340 4440 870 4566
rect 340 4374 352 4440
rect 858 4374 870 4440
rect 340 4248 870 4374
rect 340 4182 352 4248
rect 858 4182 870 4248
rect 340 4056 870 4182
rect 340 3990 352 4056
rect 858 3990 870 4056
rect 340 3864 870 3990
rect 340 3798 352 3864
rect 858 3798 870 3864
rect 340 3672 870 3798
rect 340 3606 352 3672
rect 858 3606 870 3672
rect 340 3480 870 3606
rect 340 3414 352 3480
rect 858 3414 870 3480
rect 340 3288 870 3414
rect 340 3222 352 3288
rect 858 3222 870 3288
rect 340 3096 870 3222
rect 340 3030 352 3096
rect 858 3030 870 3096
rect 340 2904 870 3030
rect 340 2838 352 2904
rect 858 2838 870 2904
rect 340 2712 870 2838
rect 340 2646 352 2712
rect 858 2646 870 2712
rect 340 2520 870 2646
rect 340 2454 352 2520
rect 858 2454 870 2520
rect 340 2328 870 2454
rect 340 2262 352 2328
rect 858 2262 870 2328
rect 340 2136 870 2262
rect 340 2070 352 2136
rect 858 2070 870 2136
rect 340 1999 870 2070
rect 970 21624 1500 23128
rect 970 21558 980 21624
rect 1490 21558 1500 21624
rect 970 21432 1500 21558
rect 970 21366 980 21432
rect 1490 21366 1500 21432
rect 970 21240 1500 21366
rect 970 21174 980 21240
rect 1490 21174 1500 21240
rect 970 21048 1500 21174
rect 970 20982 980 21048
rect 1490 20982 1500 21048
rect 970 20856 1500 20982
rect 970 20790 980 20856
rect 1490 20790 1500 20856
rect 970 20664 1500 20790
rect 970 20598 980 20664
rect 1490 20598 1500 20664
rect 970 20472 1500 20598
rect 970 20406 980 20472
rect 1490 20406 1500 20472
rect 970 20280 1500 20406
rect 970 20214 980 20280
rect 1490 20214 1500 20280
rect 970 20088 1500 20214
rect 970 20022 980 20088
rect 1490 20022 1500 20088
rect 970 19896 1500 20022
rect 970 19830 980 19896
rect 1490 19830 1500 19896
rect 970 19704 1500 19830
rect 970 19638 980 19704
rect 1490 19638 1500 19704
rect 970 19512 1500 19638
rect 970 19446 980 19512
rect 1490 19446 1500 19512
rect 970 19320 1500 19446
rect 970 19254 980 19320
rect 1490 19254 1500 19320
rect 970 19128 1500 19254
rect 970 19062 980 19128
rect 1490 19062 1500 19128
rect 970 18936 1500 19062
rect 970 18870 980 18936
rect 1490 18870 1500 18936
rect 970 18744 1500 18870
rect 970 18678 980 18744
rect 1490 18678 1500 18744
rect 970 18552 1500 18678
rect 970 18486 980 18552
rect 1490 18486 1500 18552
rect 970 18360 1500 18486
rect 970 18294 980 18360
rect 1490 18294 1500 18360
rect 970 18168 1500 18294
rect 970 18102 980 18168
rect 1490 18102 1500 18168
rect 970 17976 1500 18102
rect 970 17910 980 17976
rect 1490 17910 1500 17976
rect 970 17784 1500 17910
rect 970 17718 980 17784
rect 1490 17718 1500 17784
rect 970 17592 1500 17718
rect 970 17526 980 17592
rect 1490 17526 1500 17592
rect 970 17400 1500 17526
rect 970 17334 980 17400
rect 1490 17334 1500 17400
rect 970 17208 1500 17334
rect 970 17142 980 17208
rect 1490 17142 1500 17208
rect 970 17016 1500 17142
rect 970 16950 980 17016
rect 1490 16950 1500 17016
rect 970 16824 1500 16950
rect 970 16758 980 16824
rect 1490 16758 1500 16824
rect 970 16632 1500 16758
rect 970 16566 980 16632
rect 1490 16566 1500 16632
rect 970 16440 1500 16566
rect 970 16374 980 16440
rect 1490 16374 1500 16440
rect 970 16248 1500 16374
rect 970 16182 980 16248
rect 1490 16182 1500 16248
rect 970 16056 1500 16182
rect 970 15990 980 16056
rect 1490 15990 1500 16056
rect 970 15864 1500 15990
rect 970 15798 980 15864
rect 1490 15798 1500 15864
rect 970 15672 1500 15798
rect 970 15606 980 15672
rect 1490 15606 1500 15672
rect 970 15480 1500 15606
rect 970 15414 980 15480
rect 1490 15414 1500 15480
rect 970 15288 1500 15414
rect 970 15222 980 15288
rect 1490 15222 1500 15288
rect 970 15096 1500 15222
rect 970 15030 980 15096
rect 1490 15030 1500 15096
rect 970 14904 1500 15030
rect 970 14838 980 14904
rect 1490 14838 1500 14904
rect 970 14712 1500 14838
rect 970 14646 980 14712
rect 1490 14646 1500 14712
rect 970 14520 1500 14646
rect 970 14454 980 14520
rect 1490 14454 1500 14520
rect 970 14328 1500 14454
rect 970 14262 980 14328
rect 1490 14262 1500 14328
rect 970 14136 1500 14262
rect 970 14070 980 14136
rect 1490 14070 1500 14136
rect 970 13944 1500 14070
rect 970 13878 980 13944
rect 1490 13878 1500 13944
rect 970 13752 1500 13878
rect 970 13686 980 13752
rect 1490 13686 1500 13752
rect 970 13560 1500 13686
rect 970 13494 980 13560
rect 1490 13494 1500 13560
rect 970 13368 1500 13494
rect 970 13302 980 13368
rect 1490 13302 1500 13368
rect 970 13176 1500 13302
rect 970 13110 980 13176
rect 1490 13110 1500 13176
rect 970 12984 1500 13110
rect 970 12918 980 12984
rect 1490 12918 1500 12984
rect 970 12792 1500 12918
rect 970 12726 980 12792
rect 1490 12726 1500 12792
rect 970 12600 1500 12726
rect 970 12534 980 12600
rect 1490 12534 1500 12600
rect 970 12408 1500 12534
rect 970 12342 980 12408
rect 1490 12342 1500 12408
rect 970 12216 1500 12342
rect 970 12150 980 12216
rect 1490 12150 1500 12216
rect 970 12024 1500 12150
rect 970 11958 980 12024
rect 1490 11958 1500 12024
rect 970 11832 1500 11958
rect 970 11766 980 11832
rect 1490 11766 1500 11832
rect 970 11640 1500 11766
rect 970 11574 980 11640
rect 1490 11574 1500 11640
rect 970 11448 1500 11574
rect 970 11382 980 11448
rect 1490 11382 1500 11448
rect 970 11256 1500 11382
rect 970 11190 980 11256
rect 1490 11190 1500 11256
rect 970 11064 1500 11190
rect 970 10998 980 11064
rect 1490 10998 1500 11064
rect 970 10872 1500 10998
rect 970 10806 980 10872
rect 1490 10806 1500 10872
rect 970 10680 1500 10806
rect 970 10614 980 10680
rect 1490 10614 1500 10680
rect 970 10488 1500 10614
rect 970 10422 980 10488
rect 1490 10422 1500 10488
rect 970 10296 1500 10422
rect 970 10230 980 10296
rect 1490 10230 1500 10296
rect 970 10104 1500 10230
rect 970 10038 980 10104
rect 1490 10038 1500 10104
rect 970 9912 1500 10038
rect 970 9846 980 9912
rect 1490 9846 1500 9912
rect 970 9720 1500 9846
rect 970 9654 980 9720
rect 1490 9654 1500 9720
rect 970 9528 1500 9654
rect 970 9462 980 9528
rect 1490 9462 1500 9528
rect 970 9336 1500 9462
rect 970 9270 980 9336
rect 1490 9270 1500 9336
rect 970 9144 1500 9270
rect 970 9078 980 9144
rect 1490 9078 1500 9144
rect 970 8952 1500 9078
rect 970 8886 980 8952
rect 1490 8886 1500 8952
rect 970 8760 1500 8886
rect 970 8694 980 8760
rect 1490 8694 1500 8760
rect 970 8568 1500 8694
rect 970 8502 980 8568
rect 1490 8502 1500 8568
rect 970 8376 1500 8502
rect 970 8310 980 8376
rect 1490 8310 1500 8376
rect 970 8184 1500 8310
rect 970 8118 980 8184
rect 1490 8118 1500 8184
rect 970 7992 1500 8118
rect 970 7926 980 7992
rect 1490 7926 1500 7992
rect 970 7800 1500 7926
rect 970 7734 980 7800
rect 1490 7734 1500 7800
rect 970 7608 1500 7734
rect 970 7542 980 7608
rect 1490 7542 1500 7608
rect 970 7416 1500 7542
rect 970 7350 980 7416
rect 1490 7350 1500 7416
rect 970 7224 1500 7350
rect 970 7158 980 7224
rect 1490 7158 1500 7224
rect 970 7032 1500 7158
rect 970 6966 980 7032
rect 1490 6966 1500 7032
rect 970 6840 1500 6966
rect 970 6774 980 6840
rect 1490 6774 1500 6840
rect 970 6648 1500 6774
rect 970 6582 980 6648
rect 1490 6582 1500 6648
rect 970 6456 1500 6582
rect 970 6390 980 6456
rect 1490 6390 1500 6456
rect 970 6264 1500 6390
rect 970 6198 980 6264
rect 1490 6198 1500 6264
rect 970 6072 1500 6198
rect 970 6006 980 6072
rect 1490 6006 1500 6072
rect 970 5880 1500 6006
rect 970 5814 980 5880
rect 1490 5814 1500 5880
rect 970 5688 1500 5814
rect 970 5622 980 5688
rect 1490 5622 1500 5688
rect 970 5496 1500 5622
rect 970 5430 980 5496
rect 1490 5430 1500 5496
rect 970 5304 1500 5430
rect 970 5238 980 5304
rect 1490 5238 1500 5304
rect 970 5112 1500 5238
rect 970 5046 980 5112
rect 1490 5046 1500 5112
rect 970 4920 1500 5046
rect 970 4854 980 4920
rect 1490 4854 1500 4920
rect 970 4728 1500 4854
rect 970 4662 980 4728
rect 1490 4662 1500 4728
rect 970 4536 1500 4662
rect 970 4470 980 4536
rect 1490 4470 1500 4536
rect 970 4344 1500 4470
rect 970 4278 980 4344
rect 1490 4278 1500 4344
rect 970 4152 1500 4278
rect 970 4086 980 4152
rect 1490 4086 1500 4152
rect 970 3960 1500 4086
rect 970 3894 980 3960
rect 1490 3894 1500 3960
rect 970 3768 1500 3894
rect 970 3702 980 3768
rect 1490 3702 1500 3768
rect 970 3576 1500 3702
rect 970 3510 980 3576
rect 1490 3510 1500 3576
rect 970 3384 1500 3510
rect 970 3318 980 3384
rect 1490 3318 1500 3384
rect 970 3192 1500 3318
rect 970 3126 980 3192
rect 1490 3126 1500 3192
rect 970 3000 1500 3126
rect 970 2934 980 3000
rect 1490 2934 1500 3000
rect 970 2808 1500 2934
rect 970 2742 980 2808
rect 1490 2742 1500 2808
rect 970 2616 1500 2742
rect 970 2550 980 2616
rect 1490 2550 1500 2616
rect 970 2424 1500 2550
rect 970 2358 980 2424
rect 1490 2358 1500 2424
rect 970 2232 1500 2358
rect 970 2166 980 2232
rect 1490 2166 1500 2232
rect 970 2040 1500 2166
rect 339 1944 871 1999
rect 339 1933 352 1944
rect 340 1878 352 1933
rect 858 1933 871 1944
rect 970 1974 980 2040
rect 1490 1974 1500 2040
rect 858 1878 870 1933
rect 340 1809 870 1878
rect 970 1848 1500 1974
rect 339 1752 871 1809
rect 339 1743 352 1752
rect 340 1686 352 1743
rect 858 1743 871 1752
rect 970 1782 980 1848
rect 1490 1782 1500 1848
rect 858 1686 870 1743
rect 340 1615 870 1686
rect 970 1656 1500 1782
rect 339 1560 871 1615
rect 339 1549 352 1560
rect 340 1494 352 1549
rect 858 1549 871 1560
rect 970 1590 980 1656
rect 1490 1590 1500 1656
rect 858 1494 870 1549
rect 340 1425 870 1494
rect 970 1464 1500 1590
rect 339 1368 871 1425
rect 339 1359 352 1368
rect 340 1302 352 1359
rect 858 1359 871 1368
rect 970 1398 980 1464
rect 1490 1398 1500 1464
rect 858 1302 870 1359
rect 340 1233 870 1302
rect 970 1272 1500 1398
rect 339 1176 871 1233
rect 339 1167 352 1176
rect 340 1110 352 1167
rect 858 1167 871 1176
rect 970 1206 980 1272
rect 1490 1206 1500 1272
rect 858 1110 870 1167
rect 340 1039 870 1110
rect 970 1080 1500 1206
rect 339 984 871 1039
rect 339 973 352 984
rect 340 918 352 973
rect 858 973 871 984
rect 970 1014 980 1080
rect 1490 1014 1500 1080
rect 858 918 870 973
rect 340 849 870 918
rect 970 888 1500 1014
rect 339 792 871 849
rect 339 783 352 792
rect 340 726 352 783
rect 858 783 871 792
rect 970 822 980 888
rect 1490 822 1500 888
rect 858 726 870 783
rect 340 657 870 726
rect 970 696 1500 822
rect 339 600 871 657
rect 339 591 352 600
rect 340 534 352 591
rect 858 591 871 600
rect 970 630 980 696
rect 1490 630 1500 696
rect 858 534 870 591
rect 340 0 870 534
rect 970 0 1500 630
rect 1600 0 1840 44848
<< labels >>
rlabel metal4 0 0 240 44848 1 VGND
port 1 n ground input
rlabel metal4 1600 0 1840 44848 1 VGND
port 1 n ground input
rlabel metal4 340 0 870 44848 1 VPWR
port 2 n power input
rlabel metal4 970 0 1500 44848 1 GPWR
port 3 n power output
rlabel metal4 0 45052 1840 45152 1 ctrl
port 4 n signal input
<< end >>
