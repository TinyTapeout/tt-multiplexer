magic
tech sky130A
magscale 1 2
timestamp 1520179892
<< checkpaint >>
rect -1239 -1240 10328 16120
<< metal3 >>
rect 4501 14832 9060 14860
rect 4501 10128 4509 14832
rect 8493 10128 9060 14832
rect 4501 10060 9060 10128
rect 21 9742 9063 9770
rect 21 5198 29 9742
rect 4013 5198 9063 9742
rect 21 5108 9063 5198
rect 4501 4787 9068 4809
rect 4501 83 4509 4787
rect 8493 83 9068 4787
rect 4501 20 9068 83
<< via3 >>
rect 4509 10128 8493 14832
rect 29 5198 4013 9742
rect 4509 83 8493 4787
<< properties >>
string FIXED_BBOX 0 0 9080 14920
<< end >>
