magic
tech sky130A
magscale 1 2
timestamp 1718285629
<< metal1 >>
rect 1734 44026 1786 44032
rect 1734 98 1786 104
<< via1 >>
rect 166 44956 504 45098
rect 636 44956 1674 45098
rect 166 44688 418 44830
rect 722 44688 1674 44830
rect 32 44124 190 44596
rect 1650 44124 1808 44596
rect 1734 104 1786 44026
<< metal2 >>
rect 542 45119 598 45128
rect 160 44956 166 45098
rect 504 44956 510 45098
rect 160 44688 166 44830
rect 418 44688 424 44830
rect 630 44956 636 45098
rect 1674 44956 1680 45098
rect 542 44770 598 44779
rect 716 44688 722 44830
rect 1674 44688 1680 44830
rect 32 44596 190 44602
rect 544 44520 596 44684
rect 1650 44596 1808 44602
rect 32 44118 190 44124
rect 222 44053 274 44468
rect 990 44200 1212 44418
rect 60 43999 274 44053
rect 60 43899 192 43999
rect 994 43935 1212 44200
rect 1650 44118 1808 44124
rect 1734 44027 1790 44036
rect 60 231 138 43899
rect 1786 43878 1790 43887
rect 1734 98 1786 104
<< via2 >>
rect 169 44961 415 45030
rect 169 44756 415 44825
rect 542 44779 598 45119
rect 725 44961 1671 45030
rect 725 44756 1671 44825
rect 115 44127 185 44593
rect 1655 44127 1724 44593
rect 1734 44026 1790 44027
rect 1734 43887 1786 44026
rect 1786 43887 1790 44026
<< metal3 >>
rect 535 45146 605 45152
rect 110 45030 424 45035
rect 110 44961 169 45030
rect 415 44961 424 45030
rect 110 44956 424 44961
rect 110 44842 190 44956
rect 110 44124 111 44842
rect 189 44830 190 44842
rect 535 44954 536 45146
rect 604 44954 605 45146
rect 189 44825 424 44830
rect 415 44756 424 44825
rect 535 44779 542 44954
rect 598 44779 605 44954
rect 535 44770 605 44779
rect 716 45030 1680 45035
rect 716 44961 725 45030
rect 1671 44961 1680 45030
rect 716 44956 1680 44961
rect 716 44848 795 44956
rect 716 44847 1045 44848
rect 189 44751 424 44756
rect 189 44519 190 44751
rect 716 44689 722 44847
rect 1039 44830 1045 44847
rect 1039 44825 1680 44830
rect 1671 44756 1680 44825
rect 1039 44751 1680 44756
rect 1039 44689 1045 44751
rect 716 44688 1045 44689
rect 1650 44593 1729 44602
rect 1650 44519 1655 44593
rect 189 44440 1655 44519
rect 189 44124 190 44440
rect 110 44118 190 44124
rect 1650 44127 1655 44440
rect 1724 44127 1729 44593
rect 1650 44118 1729 44127
rect 822 44031 1795 44032
rect 822 43883 828 44031
rect 1034 44027 1795 44031
rect 1034 43887 1734 44027
rect 1790 43887 1795 44027
rect 1034 43883 1795 43887
rect 822 43882 1795 43883
<< via3 >>
rect 111 44825 189 44842
rect 536 45119 604 45146
rect 536 44954 542 45119
rect 542 44954 598 45119
rect 598 44954 604 45119
rect 111 44756 169 44825
rect 169 44756 189 44825
rect 111 44593 189 44756
rect 111 44127 115 44593
rect 115 44127 185 44593
rect 185 44127 189 44593
rect 722 44825 1039 44847
rect 722 44756 725 44825
rect 725 44756 1039 44825
rect 722 44689 1039 44756
rect 111 44124 189 44127
rect 828 43883 1034 44031
<< metal4 >>
rect 0 45146 1840 45152
rect 0 45052 536 45146
rect 535 44954 536 45052
rect 604 45052 1840 45146
rect 604 44954 605 45052
rect 535 44948 605 44954
rect 0 44842 240 44848
rect 0 44124 111 44842
rect 189 44124 240 44842
rect 0 0 240 44124
rect 340 44847 1040 44848
rect 340 44689 722 44847
rect 1039 44689 1040 44847
rect 340 44031 1040 44689
rect 340 43883 828 44031
rect 1034 43883 1040 44031
rect 340 0 1040 43883
rect 1140 0 1840 44848
use cap_gpwr  cap_gpwr_0
timestamp 1718097123
transform 1 0 0 0 1 3440
box 0 0 1840 4000
use cap_gpwr  cap_gpwr_1
timestamp 1718097123
transform 1 0 0 0 1 37712
box 0 0 1840 4000
use cap_gpwr  cap_gpwr_2
timestamp 1718097123
transform 1 0 0 0 1 14864
box 0 0 1840 4000
use cap_gpwr  cap_gpwr_3
timestamp 1718097123
transform 1 0 0 0 1 26288
box 0 0 1840 4000
use cap_vpwr  cap_vpwr_0
timestamp 1718097035
transform 1 0 0 0 1 9152
box 0 0 1840 4000
use cap_vpwr  cap_vpwr_1
timestamp 1718097035
transform 1 0 0 0 1 32000
box 0 0 1840 4000
use ckt  ckt_0
timestamp 1718271279
transform 1 0 0 0 1 608
box 0 0 1840 1120
use ckt  ckt_1
timestamp 1718271279
transform 1 0 0 0 1 2024
box 0 0 1840 1120
use ckt  ckt_2
timestamp 1718271279
transform 1 0 0 0 1 7736
box 0 0 1840 1120
use ckt  ckt_3
timestamp 1718271279
transform 1 0 0 0 1 13448
box 0 0 1840 1120
use ckt  ckt_4
timestamp 1718271279
transform 1 0 0 0 1 19576
box 0 0 1840 1120
use ckt  ckt_5
timestamp 1718271279
transform 1 0 0 0 1 20796
box 0 0 1840 1120
use ckt  ckt_6
timestamp 1718271279
transform 1 0 0 0 1 22016
box 0 0 1840 1120
use ckt  ckt_7
timestamp 1718271279
transform 1 0 0 0 1 23236
box 0 0 1840 1120
use ckt  ckt_8
timestamp 1718271279
transform 1 0 0 0 1 24456
box 0 0 1840 1120
use ckt  ckt_9
timestamp 1718271279
transform 1 0 0 0 1 30584
box 0 0 1840 1120
use ckt  ckt_10
timestamp 1718271279
transform 1 0 0 0 1 36296
box 0 0 1840 1120
use ckt  ckt_11
timestamp 1718271279
transform 1 0 0 0 1 42008
box 0 0 1840 1120
use discharge  discharge_0
timestamp 1718199492
transform 1 0 0 0 -1 44622
box 12 0 1828 524
use gate_inv  gate_inv_0
timestamp 1718283393
transform 1 0 0 0 -1 45128
box 13 0 1827 470
use pwr_pmos  pwr_pmos_0
timestamp 1718204978
transform -1 0 1810 0 1 68
box 0 0 1780 43994
<< labels >>
flabel metal4 s 0 0 240 44848 0 FreeSans 320 0 0 0 VGND
port 1 nsew ground input
flabel metal4 s 340 0 1040 44848 0 FreeSans 320 0 0 0 VPWR
port 2 nsew power input
flabel metal4 s 1140 0 1840 44848 0 FreeSans 320 0 0 0 GPWR
port 3 nsew power output
flabel metal4 s 0 45052 1840 45152 0 FreeSans 320 0 0 0 ctrl
port 4 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 1840 45152
<< end >>
