magic
tech sky130A
timestamp 1718532220
<< pwell >>
rect 0 0 836 282
<< mvnmos >>
rect 138 102 238 202
rect 278 102 378 202
rect 458 102 558 202
rect 598 102 698 202
<< mvndiff >>
rect 386 211 450 215
rect 386 202 392 211
rect 67 198 138 202
rect 67 106 73 198
rect 124 106 138 198
rect 67 102 138 106
rect 238 102 278 202
rect 378 106 392 202
rect 444 202 450 211
rect 444 106 458 202
rect 378 102 458 106
rect 558 102 598 202
rect 698 198 769 202
rect 698 106 712 198
rect 763 106 769 198
rect 698 102 769 106
<< mvndiffc >>
rect 73 106 124 198
rect 392 106 444 211
rect 712 106 763 198
<< mvpsubdiff >>
rect 13 252 45 269
rect 791 252 823 269
rect 13 237 30 252
rect 806 237 823 252
rect 13 30 30 45
rect 806 30 823 45
rect 13 13 45 30
rect 791 13 823 30
<< mvpsubdiffcont >>
rect 45 252 791 269
rect 13 45 30 237
rect 806 45 823 237
rect 45 13 791 30
<< poly >>
rect 138 202 238 215
rect 278 202 378 215
rect 458 202 558 215
rect 598 202 698 215
rect 138 86 238 102
rect 278 86 378 102
rect 458 86 558 102
rect 598 86 698 102
rect 138 81 698 86
rect 138 64 157 81
rect 679 64 698 81
rect 138 59 698 64
<< polycont >>
rect 157 64 679 81
<< locali >>
rect 13 252 45 269
rect 791 252 823 269
rect 13 237 30 252
rect 806 237 823 252
rect 386 216 450 219
rect 386 105 389 216
rect 447 105 450 216
rect 386 98 450 105
rect 149 64 157 81
rect 679 64 687 81
rect 13 30 30 45
rect 806 30 823 45
rect 13 13 45 30
rect 791 13 823 30
<< viali >>
rect 45 252 791 269
rect 13 45 30 237
rect 67 198 130 206
rect 67 106 73 198
rect 73 106 124 198
rect 124 106 130 198
rect 67 98 130 106
rect 389 211 447 216
rect 389 106 392 211
rect 392 106 444 211
rect 444 106 447 211
rect 389 105 447 106
rect 706 198 769 206
rect 706 106 712 198
rect 712 106 763 198
rect 763 106 769 198
rect 706 98 769 106
rect 157 64 679 81
rect 806 45 823 237
rect 45 13 791 30
<< metal1 >>
rect 10 269 826 272
rect 10 252 45 269
rect 791 252 826 269
rect 10 249 826 252
rect 10 237 133 249
rect 10 45 13 237
rect 30 206 133 237
rect 703 237 826 249
rect 30 98 67 206
rect 130 98 133 206
rect 383 112 386 221
rect 450 112 453 221
rect 383 105 389 112
rect 447 105 453 112
rect 383 102 453 105
rect 703 206 806 237
rect 30 45 133 98
rect 703 98 706 206
rect 769 98 806 206
rect 149 61 152 87
rect 362 84 365 87
rect 471 84 474 87
rect 362 81 474 84
rect 362 61 474 64
rect 684 61 687 87
rect 10 33 133 45
rect 703 45 806 98
rect 823 45 826 237
rect 703 33 826 45
rect 10 30 826 33
rect 10 13 45 30
rect 791 13 826 30
rect 10 10 826 13
<< via1 >>
rect 386 216 450 221
rect 386 112 389 216
rect 389 112 447 216
rect 447 112 450 216
rect 152 81 362 87
rect 474 81 684 87
rect 152 64 157 81
rect 157 64 362 81
rect 474 64 679 81
rect 679 64 684 81
rect 152 61 362 64
rect 474 61 684 64
<< metal2 >>
rect 383 112 386 221
rect 450 112 453 221
rect 149 61 152 87
rect 362 61 474 87
rect 684 61 687 87
<< end >>
