magic
tech sky130A
magscale 1 2
timestamp 1718087245
<< nwell >>
rect 0 0 1780 21290
<< pmos >>
rect 130 21079 1580 21109
rect 130 20993 1580 21023
rect 130 20907 1580 20937
rect 130 20821 1580 20851
rect 130 20735 1580 20765
rect 130 20649 1580 20679
rect 130 20563 1580 20593
rect 130 20477 1580 20507
rect 130 20391 1580 20421
rect 130 20305 1580 20335
rect 130 20219 1580 20249
rect 130 20133 1580 20163
rect 130 20047 1580 20077
rect 130 19961 1580 19991
rect 130 19875 1580 19905
rect 130 19789 1580 19819
rect 130 19703 1580 19733
rect 130 19617 1580 19647
rect 130 19531 1580 19561
rect 130 19445 1580 19475
rect 130 19359 1580 19389
rect 130 19273 1580 19303
rect 130 19187 1580 19217
rect 130 19101 1580 19131
rect 130 19015 1580 19045
rect 130 18929 1580 18959
rect 130 18843 1580 18873
rect 130 18757 1580 18787
rect 130 18671 1580 18701
rect 130 18585 1580 18615
rect 130 18499 1580 18529
rect 130 18413 1580 18443
rect 130 18327 1580 18357
rect 130 18241 1580 18271
rect 130 18155 1580 18185
rect 130 18069 1580 18099
rect 130 17983 1580 18013
rect 130 17897 1580 17927
rect 130 17811 1580 17841
rect 130 17725 1580 17755
rect 130 17639 1580 17669
rect 130 17553 1580 17583
rect 130 17467 1580 17497
rect 130 17381 1580 17411
rect 130 17295 1580 17325
rect 130 17209 1580 17239
rect 130 17123 1580 17153
rect 130 17037 1580 17067
rect 130 16951 1580 16981
rect 130 16865 1580 16895
rect 130 16779 1580 16809
rect 130 16693 1580 16723
rect 130 16607 1580 16637
rect 130 16521 1580 16551
rect 130 16435 1580 16465
rect 130 16349 1580 16379
rect 130 16263 1580 16293
rect 130 16177 1580 16207
rect 130 16091 1580 16121
rect 130 16005 1580 16035
rect 130 15919 1580 15949
rect 130 15833 1580 15863
rect 130 15747 1580 15777
rect 130 15661 1580 15691
rect 130 15575 1580 15605
rect 130 15489 1580 15519
rect 130 15403 1580 15433
rect 130 15317 1580 15347
rect 130 15231 1580 15261
rect 130 15145 1580 15175
rect 130 15059 1580 15089
rect 130 14973 1580 15003
rect 130 14887 1580 14917
rect 130 14801 1580 14831
rect 130 14715 1580 14745
rect 130 14629 1580 14659
rect 130 14543 1580 14573
rect 130 14457 1580 14487
rect 130 14371 1580 14401
rect 130 14285 1580 14315
rect 130 14199 1580 14229
rect 130 14113 1580 14143
rect 130 14027 1580 14057
rect 130 13941 1580 13971
rect 130 13855 1580 13885
rect 130 13769 1580 13799
rect 130 13683 1580 13713
rect 130 13597 1580 13627
rect 130 13511 1580 13541
rect 130 13425 1580 13455
rect 130 13339 1580 13369
rect 130 13253 1580 13283
rect 130 13167 1580 13197
rect 130 13081 1580 13111
rect 130 12995 1580 13025
rect 130 12909 1580 12939
rect 130 12823 1580 12853
rect 130 12737 1580 12767
rect 130 12651 1580 12681
rect 130 12565 1580 12595
rect 130 12479 1580 12509
rect 130 12393 1580 12423
rect 130 12307 1580 12337
rect 130 12221 1580 12251
rect 130 12135 1580 12165
rect 130 12049 1580 12079
rect 130 11963 1580 11993
rect 130 11877 1580 11907
rect 130 11791 1580 11821
rect 130 11705 1580 11735
rect 130 11619 1580 11649
rect 130 11533 1580 11563
rect 130 11447 1580 11477
rect 130 11361 1580 11391
rect 130 11275 1580 11305
rect 130 11189 1580 11219
rect 130 11103 1580 11133
rect 130 11017 1580 11047
rect 130 10931 1580 10961
rect 130 10845 1580 10875
rect 130 10759 1580 10789
rect 130 10673 1580 10703
rect 130 10587 1580 10617
rect 130 10501 1580 10531
rect 130 10415 1580 10445
rect 130 10329 1580 10359
rect 130 10243 1580 10273
rect 130 10157 1580 10187
rect 130 10071 1580 10101
rect 130 9985 1580 10015
rect 130 9899 1580 9929
rect 130 9813 1580 9843
rect 130 9727 1580 9757
rect 130 9641 1580 9671
rect 130 9555 1580 9585
rect 130 9469 1580 9499
rect 130 9383 1580 9413
rect 130 9297 1580 9327
rect 130 9211 1580 9241
rect 130 9125 1580 9155
rect 130 9039 1580 9069
rect 130 8953 1580 8983
rect 130 8867 1580 8897
rect 130 8781 1580 8811
rect 130 8695 1580 8725
rect 130 8609 1580 8639
rect 130 8523 1580 8553
rect 130 8437 1580 8467
rect 130 8351 1580 8381
rect 130 8265 1580 8295
rect 130 8179 1580 8209
rect 130 8093 1580 8123
rect 130 8007 1580 8037
rect 130 7921 1580 7951
rect 130 7835 1580 7865
rect 130 7749 1580 7779
rect 130 7663 1580 7693
rect 130 7577 1580 7607
rect 130 7491 1580 7521
rect 130 7405 1580 7435
rect 130 7319 1580 7349
rect 130 7233 1580 7263
rect 130 7147 1580 7177
rect 130 7061 1580 7091
rect 130 6975 1580 7005
rect 130 6889 1580 6919
rect 130 6803 1580 6833
rect 130 6717 1580 6747
rect 130 6631 1580 6661
rect 130 6545 1580 6575
rect 130 6459 1580 6489
rect 130 6373 1580 6403
rect 130 6287 1580 6317
rect 130 6201 1580 6231
rect 130 6115 1580 6145
rect 130 6029 1580 6059
rect 130 5943 1580 5973
rect 130 5857 1580 5887
rect 130 5771 1580 5801
rect 130 5685 1580 5715
rect 130 5599 1580 5629
rect 130 5513 1580 5543
rect 130 5427 1580 5457
rect 130 5341 1580 5371
rect 130 5255 1580 5285
rect 130 5169 1580 5199
rect 130 5083 1580 5113
rect 130 4997 1580 5027
rect 130 4911 1580 4941
rect 130 4825 1580 4855
rect 130 4739 1580 4769
rect 130 4653 1580 4683
rect 130 4567 1580 4597
rect 130 4481 1580 4511
rect 130 4395 1580 4425
rect 130 4309 1580 4339
rect 130 4223 1580 4253
rect 130 4137 1580 4167
rect 130 4051 1580 4081
rect 130 3965 1580 3995
rect 130 3879 1580 3909
rect 130 3793 1580 3823
rect 130 3707 1580 3737
rect 130 3621 1580 3651
rect 130 3535 1580 3565
rect 130 3449 1580 3479
rect 130 3363 1580 3393
rect 130 3277 1580 3307
rect 130 3191 1580 3221
rect 130 3105 1580 3135
rect 130 3019 1580 3049
rect 130 2933 1580 2963
rect 130 2847 1580 2877
rect 130 2761 1580 2791
rect 130 2675 1580 2705
rect 130 2589 1580 2619
rect 130 2503 1580 2533
rect 130 2417 1580 2447
rect 130 2331 1580 2361
rect 130 2245 1580 2275
rect 130 2159 1580 2189
rect 130 2073 1580 2103
rect 130 1987 1580 2017
rect 130 1901 1580 1931
rect 130 1815 1580 1845
rect 130 1729 1580 1759
rect 130 1643 1580 1673
rect 130 1557 1580 1587
rect 130 1471 1580 1501
rect 130 1385 1580 1415
rect 130 1299 1580 1329
rect 130 1213 1580 1243
rect 130 1127 1580 1157
rect 130 1041 1580 1071
rect 130 955 1580 985
rect 130 869 1580 899
rect 130 783 1580 813
rect 130 697 1580 727
rect 130 611 1580 641
rect 130 525 1580 555
rect 130 439 1580 469
rect 130 353 1580 383
rect 130 267 1580 297
rect 130 181 1580 211
<< pdiff >>
rect 130 21154 1580 21166
rect 130 21120 138 21154
rect 1572 21120 1580 21154
rect 130 21109 1580 21120
rect 130 21068 1580 21079
rect 130 21034 138 21068
rect 1572 21034 1580 21068
rect 130 21023 1580 21034
rect 130 20982 1580 20993
rect 130 20948 138 20982
rect 1572 20948 1580 20982
rect 130 20937 1580 20948
rect 130 20896 1580 20907
rect 130 20862 138 20896
rect 1572 20862 1580 20896
rect 130 20851 1580 20862
rect 130 20810 1580 20821
rect 130 20776 138 20810
rect 1572 20776 1580 20810
rect 130 20765 1580 20776
rect 130 20724 1580 20735
rect 130 20690 138 20724
rect 1572 20690 1580 20724
rect 130 20679 1580 20690
rect 130 20638 1580 20649
rect 130 20604 138 20638
rect 1572 20604 1580 20638
rect 130 20593 1580 20604
rect 130 20552 1580 20563
rect 130 20518 138 20552
rect 1572 20518 1580 20552
rect 130 20507 1580 20518
rect 130 20466 1580 20477
rect 130 20432 138 20466
rect 1572 20432 1580 20466
rect 130 20421 1580 20432
rect 130 20380 1580 20391
rect 130 20346 138 20380
rect 1572 20346 1580 20380
rect 130 20335 1580 20346
rect 130 20294 1580 20305
rect 130 20260 138 20294
rect 1572 20260 1580 20294
rect 130 20249 1580 20260
rect 130 20208 1580 20219
rect 130 20174 138 20208
rect 1572 20174 1580 20208
rect 130 20163 1580 20174
rect 130 20122 1580 20133
rect 130 20088 138 20122
rect 1572 20088 1580 20122
rect 130 20077 1580 20088
rect 130 20036 1580 20047
rect 130 20002 138 20036
rect 1572 20002 1580 20036
rect 130 19991 1580 20002
rect 130 19950 1580 19961
rect 130 19916 138 19950
rect 1572 19916 1580 19950
rect 130 19905 1580 19916
rect 130 19864 1580 19875
rect 130 19830 138 19864
rect 1572 19830 1580 19864
rect 130 19819 1580 19830
rect 130 19778 1580 19789
rect 130 19744 138 19778
rect 1572 19744 1580 19778
rect 130 19733 1580 19744
rect 130 19692 1580 19703
rect 130 19658 138 19692
rect 1572 19658 1580 19692
rect 130 19647 1580 19658
rect 130 19606 1580 19617
rect 130 19572 138 19606
rect 1572 19572 1580 19606
rect 130 19561 1580 19572
rect 130 19520 1580 19531
rect 130 19486 138 19520
rect 1572 19486 1580 19520
rect 130 19475 1580 19486
rect 130 19434 1580 19445
rect 130 19400 138 19434
rect 1572 19400 1580 19434
rect 130 19389 1580 19400
rect 130 19348 1580 19359
rect 130 19314 138 19348
rect 1572 19314 1580 19348
rect 130 19303 1580 19314
rect 130 19262 1580 19273
rect 130 19228 138 19262
rect 1572 19228 1580 19262
rect 130 19217 1580 19228
rect 130 19176 1580 19187
rect 130 19142 138 19176
rect 1572 19142 1580 19176
rect 130 19131 1580 19142
rect 130 19090 1580 19101
rect 130 19056 138 19090
rect 1572 19056 1580 19090
rect 130 19045 1580 19056
rect 130 19004 1580 19015
rect 130 18970 138 19004
rect 1572 18970 1580 19004
rect 130 18959 1580 18970
rect 130 18918 1580 18929
rect 130 18884 138 18918
rect 1572 18884 1580 18918
rect 130 18873 1580 18884
rect 130 18832 1580 18843
rect 130 18798 138 18832
rect 1572 18798 1580 18832
rect 130 18787 1580 18798
rect 130 18746 1580 18757
rect 130 18712 138 18746
rect 1572 18712 1580 18746
rect 130 18701 1580 18712
rect 130 18660 1580 18671
rect 130 18626 138 18660
rect 1572 18626 1580 18660
rect 130 18615 1580 18626
rect 130 18574 1580 18585
rect 130 18540 138 18574
rect 1572 18540 1580 18574
rect 130 18529 1580 18540
rect 130 18488 1580 18499
rect 130 18454 138 18488
rect 1572 18454 1580 18488
rect 130 18443 1580 18454
rect 130 18402 1580 18413
rect 130 18368 138 18402
rect 1572 18368 1580 18402
rect 130 18357 1580 18368
rect 130 18316 1580 18327
rect 130 18282 138 18316
rect 1572 18282 1580 18316
rect 130 18271 1580 18282
rect 130 18230 1580 18241
rect 130 18196 138 18230
rect 1572 18196 1580 18230
rect 130 18185 1580 18196
rect 130 18144 1580 18155
rect 130 18110 138 18144
rect 1572 18110 1580 18144
rect 130 18099 1580 18110
rect 130 18058 1580 18069
rect 130 18024 138 18058
rect 1572 18024 1580 18058
rect 130 18013 1580 18024
rect 130 17972 1580 17983
rect 130 17938 138 17972
rect 1572 17938 1580 17972
rect 130 17927 1580 17938
rect 130 17886 1580 17897
rect 130 17852 138 17886
rect 1572 17852 1580 17886
rect 130 17841 1580 17852
rect 130 17800 1580 17811
rect 130 17766 138 17800
rect 1572 17766 1580 17800
rect 130 17755 1580 17766
rect 130 17714 1580 17725
rect 130 17680 138 17714
rect 1572 17680 1580 17714
rect 130 17669 1580 17680
rect 130 17628 1580 17639
rect 130 17594 138 17628
rect 1572 17594 1580 17628
rect 130 17583 1580 17594
rect 130 17542 1580 17553
rect 130 17508 138 17542
rect 1572 17508 1580 17542
rect 130 17497 1580 17508
rect 130 17456 1580 17467
rect 130 17422 138 17456
rect 1572 17422 1580 17456
rect 130 17411 1580 17422
rect 130 17370 1580 17381
rect 130 17336 138 17370
rect 1572 17336 1580 17370
rect 130 17325 1580 17336
rect 130 17284 1580 17295
rect 130 17250 138 17284
rect 1572 17250 1580 17284
rect 130 17239 1580 17250
rect 130 17198 1580 17209
rect 130 17164 138 17198
rect 1572 17164 1580 17198
rect 130 17153 1580 17164
rect 130 17112 1580 17123
rect 130 17078 138 17112
rect 1572 17078 1580 17112
rect 130 17067 1580 17078
rect 130 17026 1580 17037
rect 130 16992 138 17026
rect 1572 16992 1580 17026
rect 130 16981 1580 16992
rect 130 16940 1580 16951
rect 130 16906 138 16940
rect 1572 16906 1580 16940
rect 130 16895 1580 16906
rect 130 16854 1580 16865
rect 130 16820 138 16854
rect 1572 16820 1580 16854
rect 130 16809 1580 16820
rect 130 16768 1580 16779
rect 130 16734 138 16768
rect 1572 16734 1580 16768
rect 130 16723 1580 16734
rect 130 16682 1580 16693
rect 130 16648 138 16682
rect 1572 16648 1580 16682
rect 130 16637 1580 16648
rect 130 16596 1580 16607
rect 130 16562 138 16596
rect 1572 16562 1580 16596
rect 130 16551 1580 16562
rect 130 16510 1580 16521
rect 130 16476 138 16510
rect 1572 16476 1580 16510
rect 130 16465 1580 16476
rect 130 16424 1580 16435
rect 130 16390 138 16424
rect 1572 16390 1580 16424
rect 130 16379 1580 16390
rect 130 16338 1580 16349
rect 130 16304 138 16338
rect 1572 16304 1580 16338
rect 130 16293 1580 16304
rect 130 16252 1580 16263
rect 130 16218 138 16252
rect 1572 16218 1580 16252
rect 130 16207 1580 16218
rect 130 16166 1580 16177
rect 130 16132 138 16166
rect 1572 16132 1580 16166
rect 130 16121 1580 16132
rect 130 16080 1580 16091
rect 130 16046 138 16080
rect 1572 16046 1580 16080
rect 130 16035 1580 16046
rect 130 15994 1580 16005
rect 130 15960 138 15994
rect 1572 15960 1580 15994
rect 130 15949 1580 15960
rect 130 15908 1580 15919
rect 130 15874 138 15908
rect 1572 15874 1580 15908
rect 130 15863 1580 15874
rect 130 15822 1580 15833
rect 130 15788 138 15822
rect 1572 15788 1580 15822
rect 130 15777 1580 15788
rect 130 15736 1580 15747
rect 130 15702 138 15736
rect 1572 15702 1580 15736
rect 130 15691 1580 15702
rect 130 15650 1580 15661
rect 130 15616 138 15650
rect 1572 15616 1580 15650
rect 130 15605 1580 15616
rect 130 15564 1580 15575
rect 130 15530 138 15564
rect 1572 15530 1580 15564
rect 130 15519 1580 15530
rect 130 15478 1580 15489
rect 130 15444 138 15478
rect 1572 15444 1580 15478
rect 130 15433 1580 15444
rect 130 15392 1580 15403
rect 130 15358 138 15392
rect 1572 15358 1580 15392
rect 130 15347 1580 15358
rect 130 15306 1580 15317
rect 130 15272 138 15306
rect 1572 15272 1580 15306
rect 130 15261 1580 15272
rect 130 15220 1580 15231
rect 130 15186 138 15220
rect 1572 15186 1580 15220
rect 130 15175 1580 15186
rect 130 15134 1580 15145
rect 130 15100 138 15134
rect 1572 15100 1580 15134
rect 130 15089 1580 15100
rect 130 15048 1580 15059
rect 130 15014 138 15048
rect 1572 15014 1580 15048
rect 130 15003 1580 15014
rect 130 14962 1580 14973
rect 130 14928 138 14962
rect 1572 14928 1580 14962
rect 130 14917 1580 14928
rect 130 14876 1580 14887
rect 130 14842 138 14876
rect 1572 14842 1580 14876
rect 130 14831 1580 14842
rect 130 14790 1580 14801
rect 130 14756 138 14790
rect 1572 14756 1580 14790
rect 130 14745 1580 14756
rect 130 14704 1580 14715
rect 130 14670 138 14704
rect 1572 14670 1580 14704
rect 130 14659 1580 14670
rect 130 14618 1580 14629
rect 130 14584 138 14618
rect 1572 14584 1580 14618
rect 130 14573 1580 14584
rect 130 14532 1580 14543
rect 130 14498 138 14532
rect 1572 14498 1580 14532
rect 130 14487 1580 14498
rect 130 14446 1580 14457
rect 130 14412 138 14446
rect 1572 14412 1580 14446
rect 130 14401 1580 14412
rect 130 14360 1580 14371
rect 130 14326 138 14360
rect 1572 14326 1580 14360
rect 130 14315 1580 14326
rect 130 14274 1580 14285
rect 130 14240 138 14274
rect 1572 14240 1580 14274
rect 130 14229 1580 14240
rect 130 14188 1580 14199
rect 130 14154 138 14188
rect 1572 14154 1580 14188
rect 130 14143 1580 14154
rect 130 14102 1580 14113
rect 130 14068 138 14102
rect 1572 14068 1580 14102
rect 130 14057 1580 14068
rect 130 14016 1580 14027
rect 130 13982 138 14016
rect 1572 13982 1580 14016
rect 130 13971 1580 13982
rect 130 13930 1580 13941
rect 130 13896 138 13930
rect 1572 13896 1580 13930
rect 130 13885 1580 13896
rect 130 13844 1580 13855
rect 130 13810 138 13844
rect 1572 13810 1580 13844
rect 130 13799 1580 13810
rect 130 13758 1580 13769
rect 130 13724 138 13758
rect 1572 13724 1580 13758
rect 130 13713 1580 13724
rect 130 13672 1580 13683
rect 130 13638 138 13672
rect 1572 13638 1580 13672
rect 130 13627 1580 13638
rect 130 13586 1580 13597
rect 130 13552 138 13586
rect 1572 13552 1580 13586
rect 130 13541 1580 13552
rect 130 13500 1580 13511
rect 130 13466 138 13500
rect 1572 13466 1580 13500
rect 130 13455 1580 13466
rect 130 13414 1580 13425
rect 130 13380 138 13414
rect 1572 13380 1580 13414
rect 130 13369 1580 13380
rect 130 13328 1580 13339
rect 130 13294 138 13328
rect 1572 13294 1580 13328
rect 130 13283 1580 13294
rect 130 13242 1580 13253
rect 130 13208 138 13242
rect 1572 13208 1580 13242
rect 130 13197 1580 13208
rect 130 13156 1580 13167
rect 130 13122 138 13156
rect 1572 13122 1580 13156
rect 130 13111 1580 13122
rect 130 13070 1580 13081
rect 130 13036 138 13070
rect 1572 13036 1580 13070
rect 130 13025 1580 13036
rect 130 12984 1580 12995
rect 130 12950 138 12984
rect 1572 12950 1580 12984
rect 130 12939 1580 12950
rect 130 12898 1580 12909
rect 130 12864 138 12898
rect 1572 12864 1580 12898
rect 130 12853 1580 12864
rect 130 12812 1580 12823
rect 130 12778 138 12812
rect 1572 12778 1580 12812
rect 130 12767 1580 12778
rect 130 12726 1580 12737
rect 130 12692 138 12726
rect 1572 12692 1580 12726
rect 130 12681 1580 12692
rect 130 12640 1580 12651
rect 130 12606 138 12640
rect 1572 12606 1580 12640
rect 130 12595 1580 12606
rect 130 12554 1580 12565
rect 130 12520 138 12554
rect 1572 12520 1580 12554
rect 130 12509 1580 12520
rect 130 12468 1580 12479
rect 130 12434 138 12468
rect 1572 12434 1580 12468
rect 130 12423 1580 12434
rect 130 12382 1580 12393
rect 130 12348 138 12382
rect 1572 12348 1580 12382
rect 130 12337 1580 12348
rect 130 12296 1580 12307
rect 130 12262 138 12296
rect 1572 12262 1580 12296
rect 130 12251 1580 12262
rect 130 12210 1580 12221
rect 130 12176 138 12210
rect 1572 12176 1580 12210
rect 130 12165 1580 12176
rect 130 12124 1580 12135
rect 130 12090 138 12124
rect 1572 12090 1580 12124
rect 130 12079 1580 12090
rect 130 12038 1580 12049
rect 130 12004 138 12038
rect 1572 12004 1580 12038
rect 130 11993 1580 12004
rect 130 11952 1580 11963
rect 130 11918 138 11952
rect 1572 11918 1580 11952
rect 130 11907 1580 11918
rect 130 11866 1580 11877
rect 130 11832 138 11866
rect 1572 11832 1580 11866
rect 130 11821 1580 11832
rect 130 11780 1580 11791
rect 130 11746 138 11780
rect 1572 11746 1580 11780
rect 130 11735 1580 11746
rect 130 11694 1580 11705
rect 130 11660 138 11694
rect 1572 11660 1580 11694
rect 130 11649 1580 11660
rect 130 11608 1580 11619
rect 130 11574 138 11608
rect 1572 11574 1580 11608
rect 130 11563 1580 11574
rect 130 11522 1580 11533
rect 130 11488 138 11522
rect 1572 11488 1580 11522
rect 130 11477 1580 11488
rect 130 11436 1580 11447
rect 130 11402 138 11436
rect 1572 11402 1580 11436
rect 130 11391 1580 11402
rect 130 11350 1580 11361
rect 130 11316 138 11350
rect 1572 11316 1580 11350
rect 130 11305 1580 11316
rect 130 11264 1580 11275
rect 130 11230 138 11264
rect 1572 11230 1580 11264
rect 130 11219 1580 11230
rect 130 11178 1580 11189
rect 130 11144 138 11178
rect 1572 11144 1580 11178
rect 130 11133 1580 11144
rect 130 11092 1580 11103
rect 130 11058 138 11092
rect 1572 11058 1580 11092
rect 130 11047 1580 11058
rect 130 11006 1580 11017
rect 130 10972 138 11006
rect 1572 10972 1580 11006
rect 130 10961 1580 10972
rect 130 10920 1580 10931
rect 130 10886 138 10920
rect 1572 10886 1580 10920
rect 130 10875 1580 10886
rect 130 10834 1580 10845
rect 130 10800 138 10834
rect 1572 10800 1580 10834
rect 130 10789 1580 10800
rect 130 10748 1580 10759
rect 130 10714 138 10748
rect 1572 10714 1580 10748
rect 130 10703 1580 10714
rect 130 10662 1580 10673
rect 130 10628 138 10662
rect 1572 10628 1580 10662
rect 130 10617 1580 10628
rect 130 10576 1580 10587
rect 130 10542 138 10576
rect 1572 10542 1580 10576
rect 130 10531 1580 10542
rect 130 10490 1580 10501
rect 130 10456 138 10490
rect 1572 10456 1580 10490
rect 130 10445 1580 10456
rect 130 10404 1580 10415
rect 130 10370 138 10404
rect 1572 10370 1580 10404
rect 130 10359 1580 10370
rect 130 10318 1580 10329
rect 130 10284 138 10318
rect 1572 10284 1580 10318
rect 130 10273 1580 10284
rect 130 10232 1580 10243
rect 130 10198 138 10232
rect 1572 10198 1580 10232
rect 130 10187 1580 10198
rect 130 10146 1580 10157
rect 130 10112 138 10146
rect 1572 10112 1580 10146
rect 130 10101 1580 10112
rect 130 10060 1580 10071
rect 130 10026 138 10060
rect 1572 10026 1580 10060
rect 130 10015 1580 10026
rect 130 9974 1580 9985
rect 130 9940 138 9974
rect 1572 9940 1580 9974
rect 130 9929 1580 9940
rect 130 9888 1580 9899
rect 130 9854 138 9888
rect 1572 9854 1580 9888
rect 130 9843 1580 9854
rect 130 9802 1580 9813
rect 130 9768 138 9802
rect 1572 9768 1580 9802
rect 130 9757 1580 9768
rect 130 9716 1580 9727
rect 130 9682 138 9716
rect 1572 9682 1580 9716
rect 130 9671 1580 9682
rect 130 9630 1580 9641
rect 130 9596 138 9630
rect 1572 9596 1580 9630
rect 130 9585 1580 9596
rect 130 9544 1580 9555
rect 130 9510 138 9544
rect 1572 9510 1580 9544
rect 130 9499 1580 9510
rect 130 9458 1580 9469
rect 130 9424 138 9458
rect 1572 9424 1580 9458
rect 130 9413 1580 9424
rect 130 9372 1580 9383
rect 130 9338 138 9372
rect 1572 9338 1580 9372
rect 130 9327 1580 9338
rect 130 9286 1580 9297
rect 130 9252 138 9286
rect 1572 9252 1580 9286
rect 130 9241 1580 9252
rect 130 9200 1580 9211
rect 130 9166 138 9200
rect 1572 9166 1580 9200
rect 130 9155 1580 9166
rect 130 9114 1580 9125
rect 130 9080 138 9114
rect 1572 9080 1580 9114
rect 130 9069 1580 9080
rect 130 9028 1580 9039
rect 130 8994 138 9028
rect 1572 8994 1580 9028
rect 130 8983 1580 8994
rect 130 8942 1580 8953
rect 130 8908 138 8942
rect 1572 8908 1580 8942
rect 130 8897 1580 8908
rect 130 8856 1580 8867
rect 130 8822 138 8856
rect 1572 8822 1580 8856
rect 130 8811 1580 8822
rect 130 8770 1580 8781
rect 130 8736 138 8770
rect 1572 8736 1580 8770
rect 130 8725 1580 8736
rect 130 8684 1580 8695
rect 130 8650 138 8684
rect 1572 8650 1580 8684
rect 130 8639 1580 8650
rect 130 8598 1580 8609
rect 130 8564 138 8598
rect 1572 8564 1580 8598
rect 130 8553 1580 8564
rect 130 8512 1580 8523
rect 130 8478 138 8512
rect 1572 8478 1580 8512
rect 130 8467 1580 8478
rect 130 8426 1580 8437
rect 130 8392 138 8426
rect 1572 8392 1580 8426
rect 130 8381 1580 8392
rect 130 8340 1580 8351
rect 130 8306 138 8340
rect 1572 8306 1580 8340
rect 130 8295 1580 8306
rect 130 8254 1580 8265
rect 130 8220 138 8254
rect 1572 8220 1580 8254
rect 130 8209 1580 8220
rect 130 8168 1580 8179
rect 130 8134 138 8168
rect 1572 8134 1580 8168
rect 130 8123 1580 8134
rect 130 8082 1580 8093
rect 130 8048 138 8082
rect 1572 8048 1580 8082
rect 130 8037 1580 8048
rect 130 7996 1580 8007
rect 130 7962 138 7996
rect 1572 7962 1580 7996
rect 130 7951 1580 7962
rect 130 7910 1580 7921
rect 130 7876 138 7910
rect 1572 7876 1580 7910
rect 130 7865 1580 7876
rect 130 7824 1580 7835
rect 130 7790 138 7824
rect 1572 7790 1580 7824
rect 130 7779 1580 7790
rect 130 7738 1580 7749
rect 130 7704 138 7738
rect 1572 7704 1580 7738
rect 130 7693 1580 7704
rect 130 7652 1580 7663
rect 130 7618 138 7652
rect 1572 7618 1580 7652
rect 130 7607 1580 7618
rect 130 7566 1580 7577
rect 130 7532 138 7566
rect 1572 7532 1580 7566
rect 130 7521 1580 7532
rect 130 7480 1580 7491
rect 130 7446 138 7480
rect 1572 7446 1580 7480
rect 130 7435 1580 7446
rect 130 7394 1580 7405
rect 130 7360 138 7394
rect 1572 7360 1580 7394
rect 130 7349 1580 7360
rect 130 7308 1580 7319
rect 130 7274 138 7308
rect 1572 7274 1580 7308
rect 130 7263 1580 7274
rect 130 7222 1580 7233
rect 130 7188 138 7222
rect 1572 7188 1580 7222
rect 130 7177 1580 7188
rect 130 7136 1580 7147
rect 130 7102 138 7136
rect 1572 7102 1580 7136
rect 130 7091 1580 7102
rect 130 7050 1580 7061
rect 130 7016 138 7050
rect 1572 7016 1580 7050
rect 130 7005 1580 7016
rect 130 6964 1580 6975
rect 130 6930 138 6964
rect 1572 6930 1580 6964
rect 130 6919 1580 6930
rect 130 6878 1580 6889
rect 130 6844 138 6878
rect 1572 6844 1580 6878
rect 130 6833 1580 6844
rect 130 6792 1580 6803
rect 130 6758 138 6792
rect 1572 6758 1580 6792
rect 130 6747 1580 6758
rect 130 6706 1580 6717
rect 130 6672 138 6706
rect 1572 6672 1580 6706
rect 130 6661 1580 6672
rect 130 6620 1580 6631
rect 130 6586 138 6620
rect 1572 6586 1580 6620
rect 130 6575 1580 6586
rect 130 6534 1580 6545
rect 130 6500 138 6534
rect 1572 6500 1580 6534
rect 130 6489 1580 6500
rect 130 6448 1580 6459
rect 130 6414 138 6448
rect 1572 6414 1580 6448
rect 130 6403 1580 6414
rect 130 6362 1580 6373
rect 130 6328 138 6362
rect 1572 6328 1580 6362
rect 130 6317 1580 6328
rect 130 6276 1580 6287
rect 130 6242 138 6276
rect 1572 6242 1580 6276
rect 130 6231 1580 6242
rect 130 6190 1580 6201
rect 130 6156 138 6190
rect 1572 6156 1580 6190
rect 130 6145 1580 6156
rect 130 6104 1580 6115
rect 130 6070 138 6104
rect 1572 6070 1580 6104
rect 130 6059 1580 6070
rect 130 6018 1580 6029
rect 130 5984 138 6018
rect 1572 5984 1580 6018
rect 130 5973 1580 5984
rect 130 5932 1580 5943
rect 130 5898 138 5932
rect 1572 5898 1580 5932
rect 130 5887 1580 5898
rect 130 5846 1580 5857
rect 130 5812 138 5846
rect 1572 5812 1580 5846
rect 130 5801 1580 5812
rect 130 5760 1580 5771
rect 130 5726 138 5760
rect 1572 5726 1580 5760
rect 130 5715 1580 5726
rect 130 5674 1580 5685
rect 130 5640 138 5674
rect 1572 5640 1580 5674
rect 130 5629 1580 5640
rect 130 5588 1580 5599
rect 130 5554 138 5588
rect 1572 5554 1580 5588
rect 130 5543 1580 5554
rect 130 5502 1580 5513
rect 130 5468 138 5502
rect 1572 5468 1580 5502
rect 130 5457 1580 5468
rect 130 5416 1580 5427
rect 130 5382 138 5416
rect 1572 5382 1580 5416
rect 130 5371 1580 5382
rect 130 5330 1580 5341
rect 130 5296 138 5330
rect 1572 5296 1580 5330
rect 130 5285 1580 5296
rect 130 5244 1580 5255
rect 130 5210 138 5244
rect 1572 5210 1580 5244
rect 130 5199 1580 5210
rect 130 5158 1580 5169
rect 130 5124 138 5158
rect 1572 5124 1580 5158
rect 130 5113 1580 5124
rect 130 5072 1580 5083
rect 130 5038 138 5072
rect 1572 5038 1580 5072
rect 130 5027 1580 5038
rect 130 4986 1580 4997
rect 130 4952 138 4986
rect 1572 4952 1580 4986
rect 130 4941 1580 4952
rect 130 4900 1580 4911
rect 130 4866 138 4900
rect 1572 4866 1580 4900
rect 130 4855 1580 4866
rect 130 4814 1580 4825
rect 130 4780 138 4814
rect 1572 4780 1580 4814
rect 130 4769 1580 4780
rect 130 4728 1580 4739
rect 130 4694 138 4728
rect 1572 4694 1580 4728
rect 130 4683 1580 4694
rect 130 4642 1580 4653
rect 130 4608 138 4642
rect 1572 4608 1580 4642
rect 130 4597 1580 4608
rect 130 4556 1580 4567
rect 130 4522 138 4556
rect 1572 4522 1580 4556
rect 130 4511 1580 4522
rect 130 4470 1580 4481
rect 130 4436 138 4470
rect 1572 4436 1580 4470
rect 130 4425 1580 4436
rect 130 4384 1580 4395
rect 130 4350 138 4384
rect 1572 4350 1580 4384
rect 130 4339 1580 4350
rect 130 4298 1580 4309
rect 130 4264 138 4298
rect 1572 4264 1580 4298
rect 130 4253 1580 4264
rect 130 4212 1580 4223
rect 130 4178 138 4212
rect 1572 4178 1580 4212
rect 130 4167 1580 4178
rect 130 4126 1580 4137
rect 130 4092 138 4126
rect 1572 4092 1580 4126
rect 130 4081 1580 4092
rect 130 4040 1580 4051
rect 130 4006 138 4040
rect 1572 4006 1580 4040
rect 130 3995 1580 4006
rect 130 3954 1580 3965
rect 130 3920 138 3954
rect 1572 3920 1580 3954
rect 130 3909 1580 3920
rect 130 3868 1580 3879
rect 130 3834 138 3868
rect 1572 3834 1580 3868
rect 130 3823 1580 3834
rect 130 3782 1580 3793
rect 130 3748 138 3782
rect 1572 3748 1580 3782
rect 130 3737 1580 3748
rect 130 3696 1580 3707
rect 130 3662 138 3696
rect 1572 3662 1580 3696
rect 130 3651 1580 3662
rect 130 3610 1580 3621
rect 130 3576 138 3610
rect 1572 3576 1580 3610
rect 130 3565 1580 3576
rect 130 3524 1580 3535
rect 130 3490 138 3524
rect 1572 3490 1580 3524
rect 130 3479 1580 3490
rect 130 3438 1580 3449
rect 130 3404 138 3438
rect 1572 3404 1580 3438
rect 130 3393 1580 3404
rect 130 3352 1580 3363
rect 130 3318 138 3352
rect 1572 3318 1580 3352
rect 130 3307 1580 3318
rect 130 3266 1580 3277
rect 130 3232 138 3266
rect 1572 3232 1580 3266
rect 130 3221 1580 3232
rect 130 3180 1580 3191
rect 130 3146 138 3180
rect 1572 3146 1580 3180
rect 130 3135 1580 3146
rect 130 3094 1580 3105
rect 130 3060 138 3094
rect 1572 3060 1580 3094
rect 130 3049 1580 3060
rect 130 3008 1580 3019
rect 130 2974 138 3008
rect 1572 2974 1580 3008
rect 130 2963 1580 2974
rect 130 2922 1580 2933
rect 130 2888 138 2922
rect 1572 2888 1580 2922
rect 130 2877 1580 2888
rect 130 2836 1580 2847
rect 130 2802 138 2836
rect 1572 2802 1580 2836
rect 130 2791 1580 2802
rect 130 2750 1580 2761
rect 130 2716 138 2750
rect 1572 2716 1580 2750
rect 130 2705 1580 2716
rect 130 2664 1580 2675
rect 130 2630 138 2664
rect 1572 2630 1580 2664
rect 130 2619 1580 2630
rect 130 2578 1580 2589
rect 130 2544 138 2578
rect 1572 2544 1580 2578
rect 130 2533 1580 2544
rect 130 2492 1580 2503
rect 130 2458 138 2492
rect 1572 2458 1580 2492
rect 130 2447 1580 2458
rect 130 2406 1580 2417
rect 130 2372 138 2406
rect 1572 2372 1580 2406
rect 130 2361 1580 2372
rect 130 2320 1580 2331
rect 130 2286 138 2320
rect 1572 2286 1580 2320
rect 130 2275 1580 2286
rect 130 2234 1580 2245
rect 130 2200 138 2234
rect 1572 2200 1580 2234
rect 130 2189 1580 2200
rect 130 2148 1580 2159
rect 130 2114 138 2148
rect 1572 2114 1580 2148
rect 130 2103 1580 2114
rect 130 2062 1580 2073
rect 130 2028 138 2062
rect 1572 2028 1580 2062
rect 130 2017 1580 2028
rect 130 1976 1580 1987
rect 130 1942 138 1976
rect 1572 1942 1580 1976
rect 130 1931 1580 1942
rect 130 1890 1580 1901
rect 130 1856 138 1890
rect 1572 1856 1580 1890
rect 130 1845 1580 1856
rect 130 1804 1580 1815
rect 130 1770 138 1804
rect 1572 1770 1580 1804
rect 130 1759 1580 1770
rect 130 1718 1580 1729
rect 130 1684 138 1718
rect 1572 1684 1580 1718
rect 130 1673 1580 1684
rect 130 1632 1580 1643
rect 130 1598 138 1632
rect 1572 1598 1580 1632
rect 130 1587 1580 1598
rect 130 1546 1580 1557
rect 130 1512 138 1546
rect 1572 1512 1580 1546
rect 130 1501 1580 1512
rect 130 1460 1580 1471
rect 130 1426 138 1460
rect 1572 1426 1580 1460
rect 130 1415 1580 1426
rect 130 1374 1580 1385
rect 130 1340 138 1374
rect 1572 1340 1580 1374
rect 130 1329 1580 1340
rect 130 1288 1580 1299
rect 130 1254 138 1288
rect 1572 1254 1580 1288
rect 130 1243 1580 1254
rect 130 1202 1580 1213
rect 130 1168 138 1202
rect 1572 1168 1580 1202
rect 130 1157 1580 1168
rect 130 1116 1580 1127
rect 130 1082 138 1116
rect 1572 1082 1580 1116
rect 130 1071 1580 1082
rect 130 1030 1580 1041
rect 130 996 138 1030
rect 1572 996 1580 1030
rect 130 985 1580 996
rect 130 944 1580 955
rect 130 910 138 944
rect 1572 910 1580 944
rect 130 899 1580 910
rect 130 858 1580 869
rect 130 824 138 858
rect 1572 824 1580 858
rect 130 813 1580 824
rect 130 772 1580 783
rect 130 738 138 772
rect 1572 738 1580 772
rect 130 727 1580 738
rect 130 686 1580 697
rect 130 652 138 686
rect 1572 652 1580 686
rect 130 641 1580 652
rect 130 600 1580 611
rect 130 566 138 600
rect 1572 566 1580 600
rect 130 555 1580 566
rect 130 514 1580 525
rect 130 480 138 514
rect 1572 480 1580 514
rect 130 469 1580 480
rect 130 428 1580 439
rect 130 394 138 428
rect 1572 394 1580 428
rect 130 383 1580 394
rect 130 342 1580 353
rect 130 308 138 342
rect 1572 308 1580 342
rect 130 297 1580 308
rect 130 256 1580 267
rect 130 222 138 256
rect 1572 222 1580 256
rect 130 211 1580 222
rect 130 170 1580 181
rect 130 136 138 170
rect 1572 136 1580 170
rect 130 124 1580 136
<< pdiffc >>
rect 138 21120 1572 21154
rect 138 21034 1572 21068
rect 138 20948 1572 20982
rect 138 20862 1572 20896
rect 138 20776 1572 20810
rect 138 20690 1572 20724
rect 138 20604 1572 20638
rect 138 20518 1572 20552
rect 138 20432 1572 20466
rect 138 20346 1572 20380
rect 138 20260 1572 20294
rect 138 20174 1572 20208
rect 138 20088 1572 20122
rect 138 20002 1572 20036
rect 138 19916 1572 19950
rect 138 19830 1572 19864
rect 138 19744 1572 19778
rect 138 19658 1572 19692
rect 138 19572 1572 19606
rect 138 19486 1572 19520
rect 138 19400 1572 19434
rect 138 19314 1572 19348
rect 138 19228 1572 19262
rect 138 19142 1572 19176
rect 138 19056 1572 19090
rect 138 18970 1572 19004
rect 138 18884 1572 18918
rect 138 18798 1572 18832
rect 138 18712 1572 18746
rect 138 18626 1572 18660
rect 138 18540 1572 18574
rect 138 18454 1572 18488
rect 138 18368 1572 18402
rect 138 18282 1572 18316
rect 138 18196 1572 18230
rect 138 18110 1572 18144
rect 138 18024 1572 18058
rect 138 17938 1572 17972
rect 138 17852 1572 17886
rect 138 17766 1572 17800
rect 138 17680 1572 17714
rect 138 17594 1572 17628
rect 138 17508 1572 17542
rect 138 17422 1572 17456
rect 138 17336 1572 17370
rect 138 17250 1572 17284
rect 138 17164 1572 17198
rect 138 17078 1572 17112
rect 138 16992 1572 17026
rect 138 16906 1572 16940
rect 138 16820 1572 16854
rect 138 16734 1572 16768
rect 138 16648 1572 16682
rect 138 16562 1572 16596
rect 138 16476 1572 16510
rect 138 16390 1572 16424
rect 138 16304 1572 16338
rect 138 16218 1572 16252
rect 138 16132 1572 16166
rect 138 16046 1572 16080
rect 138 15960 1572 15994
rect 138 15874 1572 15908
rect 138 15788 1572 15822
rect 138 15702 1572 15736
rect 138 15616 1572 15650
rect 138 15530 1572 15564
rect 138 15444 1572 15478
rect 138 15358 1572 15392
rect 138 15272 1572 15306
rect 138 15186 1572 15220
rect 138 15100 1572 15134
rect 138 15014 1572 15048
rect 138 14928 1572 14962
rect 138 14842 1572 14876
rect 138 14756 1572 14790
rect 138 14670 1572 14704
rect 138 14584 1572 14618
rect 138 14498 1572 14532
rect 138 14412 1572 14446
rect 138 14326 1572 14360
rect 138 14240 1572 14274
rect 138 14154 1572 14188
rect 138 14068 1572 14102
rect 138 13982 1572 14016
rect 138 13896 1572 13930
rect 138 13810 1572 13844
rect 138 13724 1572 13758
rect 138 13638 1572 13672
rect 138 13552 1572 13586
rect 138 13466 1572 13500
rect 138 13380 1572 13414
rect 138 13294 1572 13328
rect 138 13208 1572 13242
rect 138 13122 1572 13156
rect 138 13036 1572 13070
rect 138 12950 1572 12984
rect 138 12864 1572 12898
rect 138 12778 1572 12812
rect 138 12692 1572 12726
rect 138 12606 1572 12640
rect 138 12520 1572 12554
rect 138 12434 1572 12468
rect 138 12348 1572 12382
rect 138 12262 1572 12296
rect 138 12176 1572 12210
rect 138 12090 1572 12124
rect 138 12004 1572 12038
rect 138 11918 1572 11952
rect 138 11832 1572 11866
rect 138 11746 1572 11780
rect 138 11660 1572 11694
rect 138 11574 1572 11608
rect 138 11488 1572 11522
rect 138 11402 1572 11436
rect 138 11316 1572 11350
rect 138 11230 1572 11264
rect 138 11144 1572 11178
rect 138 11058 1572 11092
rect 138 10972 1572 11006
rect 138 10886 1572 10920
rect 138 10800 1572 10834
rect 138 10714 1572 10748
rect 138 10628 1572 10662
rect 138 10542 1572 10576
rect 138 10456 1572 10490
rect 138 10370 1572 10404
rect 138 10284 1572 10318
rect 138 10198 1572 10232
rect 138 10112 1572 10146
rect 138 10026 1572 10060
rect 138 9940 1572 9974
rect 138 9854 1572 9888
rect 138 9768 1572 9802
rect 138 9682 1572 9716
rect 138 9596 1572 9630
rect 138 9510 1572 9544
rect 138 9424 1572 9458
rect 138 9338 1572 9372
rect 138 9252 1572 9286
rect 138 9166 1572 9200
rect 138 9080 1572 9114
rect 138 8994 1572 9028
rect 138 8908 1572 8942
rect 138 8822 1572 8856
rect 138 8736 1572 8770
rect 138 8650 1572 8684
rect 138 8564 1572 8598
rect 138 8478 1572 8512
rect 138 8392 1572 8426
rect 138 8306 1572 8340
rect 138 8220 1572 8254
rect 138 8134 1572 8168
rect 138 8048 1572 8082
rect 138 7962 1572 7996
rect 138 7876 1572 7910
rect 138 7790 1572 7824
rect 138 7704 1572 7738
rect 138 7618 1572 7652
rect 138 7532 1572 7566
rect 138 7446 1572 7480
rect 138 7360 1572 7394
rect 138 7274 1572 7308
rect 138 7188 1572 7222
rect 138 7102 1572 7136
rect 138 7016 1572 7050
rect 138 6930 1572 6964
rect 138 6844 1572 6878
rect 138 6758 1572 6792
rect 138 6672 1572 6706
rect 138 6586 1572 6620
rect 138 6500 1572 6534
rect 138 6414 1572 6448
rect 138 6328 1572 6362
rect 138 6242 1572 6276
rect 138 6156 1572 6190
rect 138 6070 1572 6104
rect 138 5984 1572 6018
rect 138 5898 1572 5932
rect 138 5812 1572 5846
rect 138 5726 1572 5760
rect 138 5640 1572 5674
rect 138 5554 1572 5588
rect 138 5468 1572 5502
rect 138 5382 1572 5416
rect 138 5296 1572 5330
rect 138 5210 1572 5244
rect 138 5124 1572 5158
rect 138 5038 1572 5072
rect 138 4952 1572 4986
rect 138 4866 1572 4900
rect 138 4780 1572 4814
rect 138 4694 1572 4728
rect 138 4608 1572 4642
rect 138 4522 1572 4556
rect 138 4436 1572 4470
rect 138 4350 1572 4384
rect 138 4264 1572 4298
rect 138 4178 1572 4212
rect 138 4092 1572 4126
rect 138 4006 1572 4040
rect 138 3920 1572 3954
rect 138 3834 1572 3868
rect 138 3748 1572 3782
rect 138 3662 1572 3696
rect 138 3576 1572 3610
rect 138 3490 1572 3524
rect 138 3404 1572 3438
rect 138 3318 1572 3352
rect 138 3232 1572 3266
rect 138 3146 1572 3180
rect 138 3060 1572 3094
rect 138 2974 1572 3008
rect 138 2888 1572 2922
rect 138 2802 1572 2836
rect 138 2716 1572 2750
rect 138 2630 1572 2664
rect 138 2544 1572 2578
rect 138 2458 1572 2492
rect 138 2372 1572 2406
rect 138 2286 1572 2320
rect 138 2200 1572 2234
rect 138 2114 1572 2148
rect 138 2028 1572 2062
rect 138 1942 1572 1976
rect 138 1856 1572 1890
rect 138 1770 1572 1804
rect 138 1684 1572 1718
rect 138 1598 1572 1632
rect 138 1512 1572 1546
rect 138 1426 1572 1460
rect 138 1340 1572 1374
rect 138 1254 1572 1288
rect 138 1168 1572 1202
rect 138 1082 1572 1116
rect 138 996 1572 1030
rect 138 910 1572 944
rect 138 824 1572 858
rect 138 738 1572 772
rect 138 652 1572 686
rect 138 566 1572 600
rect 138 480 1572 514
rect 138 394 1572 428
rect 138 308 1572 342
rect 138 222 1572 256
rect 138 136 1572 170
<< nsubdiff >>
rect 36 21220 100 21254
rect 1680 21220 1744 21254
rect 36 21190 70 21220
rect 1710 21190 1744 21220
rect 36 70 70 100
rect 1710 70 1744 100
rect 36 36 100 70
rect 1680 36 1744 70
<< nsubdiffcont >>
rect 100 21220 1680 21254
rect 36 100 70 21190
rect 1710 100 1744 21190
rect 100 36 1680 70
<< poly >>
rect 1618 21111 1672 21127
rect 1618 21109 1628 21111
rect 104 21079 130 21109
rect 1580 21079 1628 21109
rect 1618 21023 1628 21079
rect 104 20993 130 21023
rect 1580 20993 1628 21023
rect 1618 20937 1628 20993
rect 104 20907 130 20937
rect 1580 20907 1628 20937
rect 1618 20851 1628 20907
rect 104 20821 130 20851
rect 1580 20821 1628 20851
rect 1618 20765 1628 20821
rect 104 20735 130 20765
rect 1580 20735 1628 20765
rect 1618 20679 1628 20735
rect 104 20649 130 20679
rect 1580 20649 1628 20679
rect 1618 20593 1628 20649
rect 104 20563 130 20593
rect 1580 20563 1628 20593
rect 1618 20507 1628 20563
rect 104 20477 130 20507
rect 1580 20477 1628 20507
rect 1618 20421 1628 20477
rect 104 20391 130 20421
rect 1580 20391 1628 20421
rect 1618 20335 1628 20391
rect 104 20305 130 20335
rect 1580 20305 1628 20335
rect 1618 20249 1628 20305
rect 104 20219 130 20249
rect 1580 20219 1628 20249
rect 1618 20163 1628 20219
rect 104 20133 130 20163
rect 1580 20133 1628 20163
rect 1618 20077 1628 20133
rect 104 20047 130 20077
rect 1580 20047 1628 20077
rect 1618 19991 1628 20047
rect 104 19961 130 19991
rect 1580 19961 1628 19991
rect 1618 19905 1628 19961
rect 104 19875 130 19905
rect 1580 19875 1628 19905
rect 1618 19819 1628 19875
rect 104 19789 130 19819
rect 1580 19789 1628 19819
rect 1618 19733 1628 19789
rect 104 19703 130 19733
rect 1580 19703 1628 19733
rect 1618 19647 1628 19703
rect 104 19617 130 19647
rect 1580 19617 1628 19647
rect 1618 19561 1628 19617
rect 104 19531 130 19561
rect 1580 19531 1628 19561
rect 1618 19475 1628 19531
rect 104 19445 130 19475
rect 1580 19445 1628 19475
rect 1618 19389 1628 19445
rect 104 19359 130 19389
rect 1580 19359 1628 19389
rect 1618 19303 1628 19359
rect 104 19273 130 19303
rect 1580 19273 1628 19303
rect 1618 19217 1628 19273
rect 104 19187 130 19217
rect 1580 19187 1628 19217
rect 1618 19131 1628 19187
rect 104 19101 130 19131
rect 1580 19101 1628 19131
rect 1618 19045 1628 19101
rect 104 19015 130 19045
rect 1580 19015 1628 19045
rect 1618 18959 1628 19015
rect 104 18929 130 18959
rect 1580 18929 1628 18959
rect 1618 18873 1628 18929
rect 104 18843 130 18873
rect 1580 18843 1628 18873
rect 1618 18787 1628 18843
rect 104 18757 130 18787
rect 1580 18757 1628 18787
rect 1618 18701 1628 18757
rect 104 18671 130 18701
rect 1580 18671 1628 18701
rect 1618 18615 1628 18671
rect 104 18585 130 18615
rect 1580 18585 1628 18615
rect 1618 18529 1628 18585
rect 104 18499 130 18529
rect 1580 18499 1628 18529
rect 1618 18443 1628 18499
rect 104 18413 130 18443
rect 1580 18413 1628 18443
rect 1618 18357 1628 18413
rect 104 18327 130 18357
rect 1580 18327 1628 18357
rect 1618 18271 1628 18327
rect 104 18241 130 18271
rect 1580 18241 1628 18271
rect 1618 18185 1628 18241
rect 104 18155 130 18185
rect 1580 18155 1628 18185
rect 1618 18099 1628 18155
rect 104 18069 130 18099
rect 1580 18069 1628 18099
rect 1618 18013 1628 18069
rect 104 17983 130 18013
rect 1580 17983 1628 18013
rect 1618 17927 1628 17983
rect 104 17897 130 17927
rect 1580 17897 1628 17927
rect 1618 17841 1628 17897
rect 104 17811 130 17841
rect 1580 17811 1628 17841
rect 1618 17755 1628 17811
rect 104 17725 130 17755
rect 1580 17725 1628 17755
rect 1618 17669 1628 17725
rect 104 17639 130 17669
rect 1580 17639 1628 17669
rect 1618 17583 1628 17639
rect 104 17553 130 17583
rect 1580 17553 1628 17583
rect 1618 17497 1628 17553
rect 104 17467 130 17497
rect 1580 17467 1628 17497
rect 1618 17411 1628 17467
rect 104 17381 130 17411
rect 1580 17381 1628 17411
rect 1618 17325 1628 17381
rect 104 17295 130 17325
rect 1580 17295 1628 17325
rect 1618 17239 1628 17295
rect 104 17209 130 17239
rect 1580 17209 1628 17239
rect 1618 17153 1628 17209
rect 104 17123 130 17153
rect 1580 17123 1628 17153
rect 1618 17067 1628 17123
rect 104 17037 130 17067
rect 1580 17037 1628 17067
rect 1618 16981 1628 17037
rect 104 16951 130 16981
rect 1580 16951 1628 16981
rect 1618 16895 1628 16951
rect 104 16865 130 16895
rect 1580 16865 1628 16895
rect 1618 16809 1628 16865
rect 104 16779 130 16809
rect 1580 16779 1628 16809
rect 1618 16723 1628 16779
rect 104 16693 130 16723
rect 1580 16693 1628 16723
rect 1618 16637 1628 16693
rect 104 16607 130 16637
rect 1580 16607 1628 16637
rect 1618 16551 1628 16607
rect 104 16521 130 16551
rect 1580 16521 1628 16551
rect 1618 16465 1628 16521
rect 104 16435 130 16465
rect 1580 16435 1628 16465
rect 1618 16379 1628 16435
rect 104 16349 130 16379
rect 1580 16349 1628 16379
rect 1618 16293 1628 16349
rect 104 16263 130 16293
rect 1580 16263 1628 16293
rect 1618 16207 1628 16263
rect 104 16177 130 16207
rect 1580 16177 1628 16207
rect 1618 16121 1628 16177
rect 104 16091 130 16121
rect 1580 16091 1628 16121
rect 1618 16035 1628 16091
rect 104 16005 130 16035
rect 1580 16005 1628 16035
rect 1618 15949 1628 16005
rect 104 15919 130 15949
rect 1580 15919 1628 15949
rect 1618 15863 1628 15919
rect 104 15833 130 15863
rect 1580 15833 1628 15863
rect 1618 15777 1628 15833
rect 104 15747 130 15777
rect 1580 15747 1628 15777
rect 1618 15691 1628 15747
rect 104 15661 130 15691
rect 1580 15661 1628 15691
rect 1618 15605 1628 15661
rect 104 15575 130 15605
rect 1580 15575 1628 15605
rect 1618 15519 1628 15575
rect 104 15489 130 15519
rect 1580 15489 1628 15519
rect 1618 15433 1628 15489
rect 104 15403 130 15433
rect 1580 15403 1628 15433
rect 1618 15347 1628 15403
rect 104 15317 130 15347
rect 1580 15317 1628 15347
rect 1618 15261 1628 15317
rect 104 15231 130 15261
rect 1580 15231 1628 15261
rect 1618 15175 1628 15231
rect 104 15145 130 15175
rect 1580 15145 1628 15175
rect 1618 15089 1628 15145
rect 104 15059 130 15089
rect 1580 15059 1628 15089
rect 1618 15003 1628 15059
rect 104 14973 130 15003
rect 1580 14973 1628 15003
rect 1618 14917 1628 14973
rect 104 14887 130 14917
rect 1580 14887 1628 14917
rect 1618 14831 1628 14887
rect 104 14801 130 14831
rect 1580 14801 1628 14831
rect 1618 14745 1628 14801
rect 104 14715 130 14745
rect 1580 14715 1628 14745
rect 1618 14659 1628 14715
rect 104 14629 130 14659
rect 1580 14629 1628 14659
rect 1618 14573 1628 14629
rect 104 14543 130 14573
rect 1580 14543 1628 14573
rect 1618 14487 1628 14543
rect 104 14457 130 14487
rect 1580 14457 1628 14487
rect 1618 14401 1628 14457
rect 104 14371 130 14401
rect 1580 14371 1628 14401
rect 1618 14315 1628 14371
rect 104 14285 130 14315
rect 1580 14285 1628 14315
rect 1618 14229 1628 14285
rect 104 14199 130 14229
rect 1580 14199 1628 14229
rect 1618 14143 1628 14199
rect 104 14113 130 14143
rect 1580 14113 1628 14143
rect 1618 14057 1628 14113
rect 104 14027 130 14057
rect 1580 14027 1628 14057
rect 1618 13971 1628 14027
rect 104 13941 130 13971
rect 1580 13941 1628 13971
rect 1618 13885 1628 13941
rect 104 13855 130 13885
rect 1580 13855 1628 13885
rect 1618 13799 1628 13855
rect 104 13769 130 13799
rect 1580 13769 1628 13799
rect 1618 13713 1628 13769
rect 104 13683 130 13713
rect 1580 13683 1628 13713
rect 1618 13627 1628 13683
rect 104 13597 130 13627
rect 1580 13597 1628 13627
rect 1618 13541 1628 13597
rect 104 13511 130 13541
rect 1580 13511 1628 13541
rect 1618 13455 1628 13511
rect 104 13425 130 13455
rect 1580 13425 1628 13455
rect 1618 13369 1628 13425
rect 104 13339 130 13369
rect 1580 13339 1628 13369
rect 1618 13283 1628 13339
rect 104 13253 130 13283
rect 1580 13253 1628 13283
rect 1618 13197 1628 13253
rect 104 13167 130 13197
rect 1580 13167 1628 13197
rect 1618 13111 1628 13167
rect 104 13081 130 13111
rect 1580 13081 1628 13111
rect 1618 13025 1628 13081
rect 104 12995 130 13025
rect 1580 12995 1628 13025
rect 1618 12939 1628 12995
rect 104 12909 130 12939
rect 1580 12909 1628 12939
rect 1618 12853 1628 12909
rect 104 12823 130 12853
rect 1580 12823 1628 12853
rect 1618 12767 1628 12823
rect 104 12737 130 12767
rect 1580 12737 1628 12767
rect 1618 12681 1628 12737
rect 104 12651 130 12681
rect 1580 12651 1628 12681
rect 1618 12595 1628 12651
rect 104 12565 130 12595
rect 1580 12565 1628 12595
rect 1618 12509 1628 12565
rect 104 12479 130 12509
rect 1580 12479 1628 12509
rect 1618 12423 1628 12479
rect 104 12393 130 12423
rect 1580 12393 1628 12423
rect 1618 12337 1628 12393
rect 104 12307 130 12337
rect 1580 12307 1628 12337
rect 1618 12251 1628 12307
rect 104 12221 130 12251
rect 1580 12221 1628 12251
rect 1618 12165 1628 12221
rect 104 12135 130 12165
rect 1580 12135 1628 12165
rect 1618 12079 1628 12135
rect 104 12049 130 12079
rect 1580 12049 1628 12079
rect 1618 11993 1628 12049
rect 104 11963 130 11993
rect 1580 11963 1628 11993
rect 1618 11907 1628 11963
rect 104 11877 130 11907
rect 1580 11877 1628 11907
rect 1618 11821 1628 11877
rect 104 11791 130 11821
rect 1580 11791 1628 11821
rect 1618 11735 1628 11791
rect 104 11705 130 11735
rect 1580 11705 1628 11735
rect 1618 11649 1628 11705
rect 104 11619 130 11649
rect 1580 11619 1628 11649
rect 1618 11563 1628 11619
rect 104 11533 130 11563
rect 1580 11533 1628 11563
rect 1618 11477 1628 11533
rect 104 11447 130 11477
rect 1580 11447 1628 11477
rect 1618 11391 1628 11447
rect 104 11361 130 11391
rect 1580 11361 1628 11391
rect 1618 11305 1628 11361
rect 104 11275 130 11305
rect 1580 11275 1628 11305
rect 1618 11219 1628 11275
rect 104 11189 130 11219
rect 1580 11189 1628 11219
rect 1618 11133 1628 11189
rect 104 11103 130 11133
rect 1580 11103 1628 11133
rect 1618 11047 1628 11103
rect 104 11017 130 11047
rect 1580 11017 1628 11047
rect 1618 10961 1628 11017
rect 104 10931 130 10961
rect 1580 10931 1628 10961
rect 1618 10875 1628 10931
rect 104 10845 130 10875
rect 1580 10845 1628 10875
rect 1618 10789 1628 10845
rect 104 10759 130 10789
rect 1580 10759 1628 10789
rect 1618 10703 1628 10759
rect 104 10673 130 10703
rect 1580 10673 1628 10703
rect 1618 10617 1628 10673
rect 104 10587 130 10617
rect 1580 10587 1628 10617
rect 1618 10531 1628 10587
rect 104 10501 130 10531
rect 1580 10501 1628 10531
rect 1618 10445 1628 10501
rect 104 10415 130 10445
rect 1580 10415 1628 10445
rect 1618 10359 1628 10415
rect 104 10329 130 10359
rect 1580 10329 1628 10359
rect 1618 10273 1628 10329
rect 104 10243 130 10273
rect 1580 10243 1628 10273
rect 1618 10187 1628 10243
rect 104 10157 130 10187
rect 1580 10157 1628 10187
rect 1618 10101 1628 10157
rect 104 10071 130 10101
rect 1580 10071 1628 10101
rect 1618 10015 1628 10071
rect 104 9985 130 10015
rect 1580 9985 1628 10015
rect 1618 9929 1628 9985
rect 104 9899 130 9929
rect 1580 9899 1628 9929
rect 1618 9843 1628 9899
rect 104 9813 130 9843
rect 1580 9813 1628 9843
rect 1618 9757 1628 9813
rect 104 9727 130 9757
rect 1580 9727 1628 9757
rect 1618 9671 1628 9727
rect 104 9641 130 9671
rect 1580 9641 1628 9671
rect 1618 9585 1628 9641
rect 104 9555 130 9585
rect 1580 9555 1628 9585
rect 1618 9499 1628 9555
rect 104 9469 130 9499
rect 1580 9469 1628 9499
rect 1618 9413 1628 9469
rect 104 9383 130 9413
rect 1580 9383 1628 9413
rect 1618 9327 1628 9383
rect 104 9297 130 9327
rect 1580 9297 1628 9327
rect 1618 9241 1628 9297
rect 104 9211 130 9241
rect 1580 9211 1628 9241
rect 1618 9155 1628 9211
rect 104 9125 130 9155
rect 1580 9125 1628 9155
rect 1618 9069 1628 9125
rect 104 9039 130 9069
rect 1580 9039 1628 9069
rect 1618 8983 1628 9039
rect 104 8953 130 8983
rect 1580 8953 1628 8983
rect 1618 8897 1628 8953
rect 104 8867 130 8897
rect 1580 8867 1628 8897
rect 1618 8811 1628 8867
rect 104 8781 130 8811
rect 1580 8781 1628 8811
rect 1618 8725 1628 8781
rect 104 8695 130 8725
rect 1580 8695 1628 8725
rect 1618 8639 1628 8695
rect 104 8609 130 8639
rect 1580 8609 1628 8639
rect 1618 8553 1628 8609
rect 104 8523 130 8553
rect 1580 8523 1628 8553
rect 1618 8467 1628 8523
rect 104 8437 130 8467
rect 1580 8437 1628 8467
rect 1618 8381 1628 8437
rect 104 8351 130 8381
rect 1580 8351 1628 8381
rect 1618 8295 1628 8351
rect 104 8265 130 8295
rect 1580 8265 1628 8295
rect 1618 8209 1628 8265
rect 104 8179 130 8209
rect 1580 8179 1628 8209
rect 1618 8123 1628 8179
rect 104 8093 130 8123
rect 1580 8093 1628 8123
rect 1618 8037 1628 8093
rect 104 8007 130 8037
rect 1580 8007 1628 8037
rect 1618 7951 1628 8007
rect 104 7921 130 7951
rect 1580 7921 1628 7951
rect 1618 7865 1628 7921
rect 104 7835 130 7865
rect 1580 7835 1628 7865
rect 1618 7779 1628 7835
rect 104 7749 130 7779
rect 1580 7749 1628 7779
rect 1618 7693 1628 7749
rect 104 7663 130 7693
rect 1580 7663 1628 7693
rect 1618 7607 1628 7663
rect 104 7577 130 7607
rect 1580 7577 1628 7607
rect 1618 7521 1628 7577
rect 104 7491 130 7521
rect 1580 7491 1628 7521
rect 1618 7435 1628 7491
rect 104 7405 130 7435
rect 1580 7405 1628 7435
rect 1618 7349 1628 7405
rect 104 7319 130 7349
rect 1580 7319 1628 7349
rect 1618 7263 1628 7319
rect 104 7233 130 7263
rect 1580 7233 1628 7263
rect 1618 7177 1628 7233
rect 104 7147 130 7177
rect 1580 7147 1628 7177
rect 1618 7091 1628 7147
rect 104 7061 130 7091
rect 1580 7061 1628 7091
rect 1618 7005 1628 7061
rect 104 6975 130 7005
rect 1580 6975 1628 7005
rect 1618 6919 1628 6975
rect 104 6889 130 6919
rect 1580 6889 1628 6919
rect 1618 6833 1628 6889
rect 104 6803 130 6833
rect 1580 6803 1628 6833
rect 1618 6747 1628 6803
rect 104 6717 130 6747
rect 1580 6717 1628 6747
rect 1618 6661 1628 6717
rect 104 6631 130 6661
rect 1580 6631 1628 6661
rect 1618 6575 1628 6631
rect 104 6545 130 6575
rect 1580 6545 1628 6575
rect 1618 6489 1628 6545
rect 104 6459 130 6489
rect 1580 6459 1628 6489
rect 1618 6403 1628 6459
rect 104 6373 130 6403
rect 1580 6373 1628 6403
rect 1618 6317 1628 6373
rect 104 6287 130 6317
rect 1580 6287 1628 6317
rect 1618 6231 1628 6287
rect 104 6201 130 6231
rect 1580 6201 1628 6231
rect 1618 6145 1628 6201
rect 104 6115 130 6145
rect 1580 6115 1628 6145
rect 1618 6059 1628 6115
rect 104 6029 130 6059
rect 1580 6029 1628 6059
rect 1618 5973 1628 6029
rect 104 5943 130 5973
rect 1580 5943 1628 5973
rect 1618 5887 1628 5943
rect 104 5857 130 5887
rect 1580 5857 1628 5887
rect 1618 5801 1628 5857
rect 104 5771 130 5801
rect 1580 5771 1628 5801
rect 1618 5715 1628 5771
rect 104 5685 130 5715
rect 1580 5685 1628 5715
rect 1618 5629 1628 5685
rect 104 5599 130 5629
rect 1580 5599 1628 5629
rect 1618 5543 1628 5599
rect 104 5513 130 5543
rect 1580 5513 1628 5543
rect 1618 5457 1628 5513
rect 104 5427 130 5457
rect 1580 5427 1628 5457
rect 1618 5371 1628 5427
rect 104 5341 130 5371
rect 1580 5341 1628 5371
rect 1618 5285 1628 5341
rect 104 5255 130 5285
rect 1580 5255 1628 5285
rect 1618 5199 1628 5255
rect 104 5169 130 5199
rect 1580 5169 1628 5199
rect 1618 5113 1628 5169
rect 104 5083 130 5113
rect 1580 5083 1628 5113
rect 1618 5027 1628 5083
rect 104 4997 130 5027
rect 1580 4997 1628 5027
rect 1618 4941 1628 4997
rect 104 4911 130 4941
rect 1580 4911 1628 4941
rect 1618 4855 1628 4911
rect 104 4825 130 4855
rect 1580 4825 1628 4855
rect 1618 4769 1628 4825
rect 104 4739 130 4769
rect 1580 4739 1628 4769
rect 1618 4683 1628 4739
rect 104 4653 130 4683
rect 1580 4653 1628 4683
rect 1618 4597 1628 4653
rect 104 4567 130 4597
rect 1580 4567 1628 4597
rect 1618 4511 1628 4567
rect 104 4481 130 4511
rect 1580 4481 1628 4511
rect 1618 4425 1628 4481
rect 104 4395 130 4425
rect 1580 4395 1628 4425
rect 1618 4339 1628 4395
rect 104 4309 130 4339
rect 1580 4309 1628 4339
rect 1618 4253 1628 4309
rect 104 4223 130 4253
rect 1580 4223 1628 4253
rect 1618 4167 1628 4223
rect 104 4137 130 4167
rect 1580 4137 1628 4167
rect 1618 4081 1628 4137
rect 104 4051 130 4081
rect 1580 4051 1628 4081
rect 1618 3995 1628 4051
rect 104 3965 130 3995
rect 1580 3965 1628 3995
rect 1618 3909 1628 3965
rect 104 3879 130 3909
rect 1580 3879 1628 3909
rect 1618 3823 1628 3879
rect 104 3793 130 3823
rect 1580 3793 1628 3823
rect 1618 3737 1628 3793
rect 104 3707 130 3737
rect 1580 3707 1628 3737
rect 1618 3651 1628 3707
rect 104 3621 130 3651
rect 1580 3621 1628 3651
rect 1618 3565 1628 3621
rect 104 3535 130 3565
rect 1580 3535 1628 3565
rect 1618 3479 1628 3535
rect 104 3449 130 3479
rect 1580 3449 1628 3479
rect 1618 3393 1628 3449
rect 104 3363 130 3393
rect 1580 3363 1628 3393
rect 1618 3307 1628 3363
rect 104 3277 130 3307
rect 1580 3277 1628 3307
rect 1618 3221 1628 3277
rect 104 3191 130 3221
rect 1580 3191 1628 3221
rect 1618 3135 1628 3191
rect 104 3105 130 3135
rect 1580 3105 1628 3135
rect 1618 3049 1628 3105
rect 104 3019 130 3049
rect 1580 3019 1628 3049
rect 1618 2963 1628 3019
rect 104 2933 130 2963
rect 1580 2933 1628 2963
rect 1618 2877 1628 2933
rect 104 2847 130 2877
rect 1580 2847 1628 2877
rect 1618 2791 1628 2847
rect 104 2761 130 2791
rect 1580 2761 1628 2791
rect 1618 2705 1628 2761
rect 104 2675 130 2705
rect 1580 2675 1628 2705
rect 1618 2619 1628 2675
rect 104 2589 130 2619
rect 1580 2589 1628 2619
rect 1618 2533 1628 2589
rect 104 2503 130 2533
rect 1580 2503 1628 2533
rect 1618 2447 1628 2503
rect 104 2417 130 2447
rect 1580 2417 1628 2447
rect 1618 2361 1628 2417
rect 104 2331 130 2361
rect 1580 2331 1628 2361
rect 1618 2275 1628 2331
rect 104 2245 130 2275
rect 1580 2245 1628 2275
rect 1618 2189 1628 2245
rect 104 2159 130 2189
rect 1580 2159 1628 2189
rect 1618 2103 1628 2159
rect 104 2073 130 2103
rect 1580 2073 1628 2103
rect 1618 2017 1628 2073
rect 104 1987 130 2017
rect 1580 1987 1628 2017
rect 1618 1931 1628 1987
rect 104 1901 130 1931
rect 1580 1901 1628 1931
rect 1618 1845 1628 1901
rect 104 1815 130 1845
rect 1580 1815 1628 1845
rect 1618 1759 1628 1815
rect 104 1729 130 1759
rect 1580 1729 1628 1759
rect 1618 1673 1628 1729
rect 104 1643 130 1673
rect 1580 1643 1628 1673
rect 1618 1587 1628 1643
rect 104 1557 130 1587
rect 1580 1557 1628 1587
rect 1618 1501 1628 1557
rect 104 1471 130 1501
rect 1580 1471 1628 1501
rect 1618 1415 1628 1471
rect 104 1385 130 1415
rect 1580 1385 1628 1415
rect 1618 1329 1628 1385
rect 104 1299 130 1329
rect 1580 1299 1628 1329
rect 1618 1243 1628 1299
rect 104 1213 130 1243
rect 1580 1213 1628 1243
rect 1618 1157 1628 1213
rect 104 1127 130 1157
rect 1580 1127 1628 1157
rect 1618 1071 1628 1127
rect 104 1041 130 1071
rect 1580 1041 1628 1071
rect 1618 985 1628 1041
rect 104 955 130 985
rect 1580 955 1628 985
rect 1618 899 1628 955
rect 104 869 130 899
rect 1580 869 1628 899
rect 1618 813 1628 869
rect 104 783 130 813
rect 1580 783 1628 813
rect 1618 727 1628 783
rect 104 697 130 727
rect 1580 697 1628 727
rect 1618 641 1628 697
rect 104 611 130 641
rect 1580 611 1628 641
rect 1618 555 1628 611
rect 104 525 130 555
rect 1580 525 1628 555
rect 1618 469 1628 525
rect 104 439 130 469
rect 1580 439 1628 469
rect 1618 383 1628 439
rect 104 353 130 383
rect 1580 353 1628 383
rect 1618 297 1628 353
rect 104 267 130 297
rect 1580 267 1628 297
rect 1618 211 1628 267
rect 104 181 130 211
rect 1580 181 1628 211
rect 1618 179 1628 181
rect 1662 179 1672 21111
rect 1618 163 1672 179
<< polycont >>
rect 1628 179 1662 21111
<< locali >>
rect 36 21220 100 21254
rect 1680 21220 1744 21254
rect 36 21190 70 21220
rect 1710 21190 1744 21220
rect 122 21120 138 21154
rect 1572 21120 1588 21154
rect 1628 21111 1662 21127
rect 122 21034 138 21068
rect 1572 21034 1588 21068
rect 122 20948 138 20982
rect 1572 20948 1588 20982
rect 122 20862 138 20896
rect 1572 20862 1588 20896
rect 122 20776 138 20810
rect 1572 20776 1588 20810
rect 122 20690 138 20724
rect 1572 20690 1588 20724
rect 122 20604 138 20638
rect 1572 20604 1588 20638
rect 122 20518 138 20552
rect 1572 20518 1588 20552
rect 122 20432 138 20466
rect 1572 20432 1588 20466
rect 122 20346 138 20380
rect 1572 20346 1588 20380
rect 122 20260 138 20294
rect 1572 20260 1588 20294
rect 122 20174 138 20208
rect 1572 20174 1588 20208
rect 122 20088 138 20122
rect 1572 20088 1588 20122
rect 122 20002 138 20036
rect 1572 20002 1588 20036
rect 122 19916 138 19950
rect 1572 19916 1588 19950
rect 122 19830 138 19864
rect 1572 19830 1588 19864
rect 122 19744 138 19778
rect 1572 19744 1588 19778
rect 122 19658 138 19692
rect 1572 19658 1588 19692
rect 122 19572 138 19606
rect 1572 19572 1588 19606
rect 122 19486 138 19520
rect 1572 19486 1588 19520
rect 122 19400 138 19434
rect 1572 19400 1588 19434
rect 122 19314 138 19348
rect 1572 19314 1588 19348
rect 122 19228 138 19262
rect 1572 19228 1588 19262
rect 122 19142 138 19176
rect 1572 19142 1588 19176
rect 122 19056 138 19090
rect 1572 19056 1588 19090
rect 122 18970 138 19004
rect 1572 18970 1588 19004
rect 122 18884 138 18918
rect 1572 18884 1588 18918
rect 122 18798 138 18832
rect 1572 18798 1588 18832
rect 122 18712 138 18746
rect 1572 18712 1588 18746
rect 122 18626 138 18660
rect 1572 18626 1588 18660
rect 122 18540 138 18574
rect 1572 18540 1588 18574
rect 122 18454 138 18488
rect 1572 18454 1588 18488
rect 122 18368 138 18402
rect 1572 18368 1588 18402
rect 122 18282 138 18316
rect 1572 18282 1588 18316
rect 122 18196 138 18230
rect 1572 18196 1588 18230
rect 122 18110 138 18144
rect 1572 18110 1588 18144
rect 122 18024 138 18058
rect 1572 18024 1588 18058
rect 122 17938 138 17972
rect 1572 17938 1588 17972
rect 122 17852 138 17886
rect 1572 17852 1588 17886
rect 122 17766 138 17800
rect 1572 17766 1588 17800
rect 122 17680 138 17714
rect 1572 17680 1588 17714
rect 122 17594 138 17628
rect 1572 17594 1588 17628
rect 122 17508 138 17542
rect 1572 17508 1588 17542
rect 122 17422 138 17456
rect 1572 17422 1588 17456
rect 122 17336 138 17370
rect 1572 17336 1588 17370
rect 122 17250 138 17284
rect 1572 17250 1588 17284
rect 122 17164 138 17198
rect 1572 17164 1588 17198
rect 122 17078 138 17112
rect 1572 17078 1588 17112
rect 122 16992 138 17026
rect 1572 16992 1588 17026
rect 122 16906 138 16940
rect 1572 16906 1588 16940
rect 122 16820 138 16854
rect 1572 16820 1588 16854
rect 122 16734 138 16768
rect 1572 16734 1588 16768
rect 122 16648 138 16682
rect 1572 16648 1588 16682
rect 122 16562 138 16596
rect 1572 16562 1588 16596
rect 122 16476 138 16510
rect 1572 16476 1588 16510
rect 122 16390 138 16424
rect 1572 16390 1588 16424
rect 122 16304 138 16338
rect 1572 16304 1588 16338
rect 122 16218 138 16252
rect 1572 16218 1588 16252
rect 122 16132 138 16166
rect 1572 16132 1588 16166
rect 122 16046 138 16080
rect 1572 16046 1588 16080
rect 122 15960 138 15994
rect 1572 15960 1588 15994
rect 122 15874 138 15908
rect 1572 15874 1588 15908
rect 122 15788 138 15822
rect 1572 15788 1588 15822
rect 122 15702 138 15736
rect 1572 15702 1588 15736
rect 122 15616 138 15650
rect 1572 15616 1588 15650
rect 122 15530 138 15564
rect 1572 15530 1588 15564
rect 122 15444 138 15478
rect 1572 15444 1588 15478
rect 122 15358 138 15392
rect 1572 15358 1588 15392
rect 122 15272 138 15306
rect 1572 15272 1588 15306
rect 122 15186 138 15220
rect 1572 15186 1588 15220
rect 122 15100 138 15134
rect 1572 15100 1588 15134
rect 122 15014 138 15048
rect 1572 15014 1588 15048
rect 122 14928 138 14962
rect 1572 14928 1588 14962
rect 122 14842 138 14876
rect 1572 14842 1588 14876
rect 122 14756 138 14790
rect 1572 14756 1588 14790
rect 122 14670 138 14704
rect 1572 14670 1588 14704
rect 122 14584 138 14618
rect 1572 14584 1588 14618
rect 122 14498 138 14532
rect 1572 14498 1588 14532
rect 122 14412 138 14446
rect 1572 14412 1588 14446
rect 122 14326 138 14360
rect 1572 14326 1588 14360
rect 122 14240 138 14274
rect 1572 14240 1588 14274
rect 122 14154 138 14188
rect 1572 14154 1588 14188
rect 122 14068 138 14102
rect 1572 14068 1588 14102
rect 122 13982 138 14016
rect 1572 13982 1588 14016
rect 122 13896 138 13930
rect 1572 13896 1588 13930
rect 122 13810 138 13844
rect 1572 13810 1588 13844
rect 122 13724 138 13758
rect 1572 13724 1588 13758
rect 122 13638 138 13672
rect 1572 13638 1588 13672
rect 122 13552 138 13586
rect 1572 13552 1588 13586
rect 122 13466 138 13500
rect 1572 13466 1588 13500
rect 122 13380 138 13414
rect 1572 13380 1588 13414
rect 122 13294 138 13328
rect 1572 13294 1588 13328
rect 122 13208 138 13242
rect 1572 13208 1588 13242
rect 122 13122 138 13156
rect 1572 13122 1588 13156
rect 122 13036 138 13070
rect 1572 13036 1588 13070
rect 122 12950 138 12984
rect 1572 12950 1588 12984
rect 122 12864 138 12898
rect 1572 12864 1588 12898
rect 122 12778 138 12812
rect 1572 12778 1588 12812
rect 122 12692 138 12726
rect 1572 12692 1588 12726
rect 122 12606 138 12640
rect 1572 12606 1588 12640
rect 122 12520 138 12554
rect 1572 12520 1588 12554
rect 122 12434 138 12468
rect 1572 12434 1588 12468
rect 122 12348 138 12382
rect 1572 12348 1588 12382
rect 122 12262 138 12296
rect 1572 12262 1588 12296
rect 122 12176 138 12210
rect 1572 12176 1588 12210
rect 122 12090 138 12124
rect 1572 12090 1588 12124
rect 122 12004 138 12038
rect 1572 12004 1588 12038
rect 122 11918 138 11952
rect 1572 11918 1588 11952
rect 122 11832 138 11866
rect 1572 11832 1588 11866
rect 122 11746 138 11780
rect 1572 11746 1588 11780
rect 122 11660 138 11694
rect 1572 11660 1588 11694
rect 122 11574 138 11608
rect 1572 11574 1588 11608
rect 122 11488 138 11522
rect 1572 11488 1588 11522
rect 122 11402 138 11436
rect 1572 11402 1588 11436
rect 122 11316 138 11350
rect 1572 11316 1588 11350
rect 122 11230 138 11264
rect 1572 11230 1588 11264
rect 122 11144 138 11178
rect 1572 11144 1588 11178
rect 122 11058 138 11092
rect 1572 11058 1588 11092
rect 122 10972 138 11006
rect 1572 10972 1588 11006
rect 122 10886 138 10920
rect 1572 10886 1588 10920
rect 122 10800 138 10834
rect 1572 10800 1588 10834
rect 122 10714 138 10748
rect 1572 10714 1588 10748
rect 122 10628 138 10662
rect 1572 10628 1588 10662
rect 122 10542 138 10576
rect 1572 10542 1588 10576
rect 122 10456 138 10490
rect 1572 10456 1588 10490
rect 122 10370 138 10404
rect 1572 10370 1588 10404
rect 122 10284 138 10318
rect 1572 10284 1588 10318
rect 122 10198 138 10232
rect 1572 10198 1588 10232
rect 122 10112 138 10146
rect 1572 10112 1588 10146
rect 122 10026 138 10060
rect 1572 10026 1588 10060
rect 122 9940 138 9974
rect 1572 9940 1588 9974
rect 122 9854 138 9888
rect 1572 9854 1588 9888
rect 122 9768 138 9802
rect 1572 9768 1588 9802
rect 122 9682 138 9716
rect 1572 9682 1588 9716
rect 122 9596 138 9630
rect 1572 9596 1588 9630
rect 122 9510 138 9544
rect 1572 9510 1588 9544
rect 122 9424 138 9458
rect 1572 9424 1588 9458
rect 122 9338 138 9372
rect 1572 9338 1588 9372
rect 122 9252 138 9286
rect 1572 9252 1588 9286
rect 122 9166 138 9200
rect 1572 9166 1588 9200
rect 122 9080 138 9114
rect 1572 9080 1588 9114
rect 122 8994 138 9028
rect 1572 8994 1588 9028
rect 122 8908 138 8942
rect 1572 8908 1588 8942
rect 122 8822 138 8856
rect 1572 8822 1588 8856
rect 122 8736 138 8770
rect 1572 8736 1588 8770
rect 122 8650 138 8684
rect 1572 8650 1588 8684
rect 122 8564 138 8598
rect 1572 8564 1588 8598
rect 122 8478 138 8512
rect 1572 8478 1588 8512
rect 122 8392 138 8426
rect 1572 8392 1588 8426
rect 122 8306 138 8340
rect 1572 8306 1588 8340
rect 122 8220 138 8254
rect 1572 8220 1588 8254
rect 122 8134 138 8168
rect 1572 8134 1588 8168
rect 122 8048 138 8082
rect 1572 8048 1588 8082
rect 122 7962 138 7996
rect 1572 7962 1588 7996
rect 122 7876 138 7910
rect 1572 7876 1588 7910
rect 122 7790 138 7824
rect 1572 7790 1588 7824
rect 122 7704 138 7738
rect 1572 7704 1588 7738
rect 122 7618 138 7652
rect 1572 7618 1588 7652
rect 122 7532 138 7566
rect 1572 7532 1588 7566
rect 122 7446 138 7480
rect 1572 7446 1588 7480
rect 122 7360 138 7394
rect 1572 7360 1588 7394
rect 122 7274 138 7308
rect 1572 7274 1588 7308
rect 122 7188 138 7222
rect 1572 7188 1588 7222
rect 122 7102 138 7136
rect 1572 7102 1588 7136
rect 122 7016 138 7050
rect 1572 7016 1588 7050
rect 122 6930 138 6964
rect 1572 6930 1588 6964
rect 122 6844 138 6878
rect 1572 6844 1588 6878
rect 122 6758 138 6792
rect 1572 6758 1588 6792
rect 122 6672 138 6706
rect 1572 6672 1588 6706
rect 122 6586 138 6620
rect 1572 6586 1588 6620
rect 122 6500 138 6534
rect 1572 6500 1588 6534
rect 122 6414 138 6448
rect 1572 6414 1588 6448
rect 122 6328 138 6362
rect 1572 6328 1588 6362
rect 122 6242 138 6276
rect 1572 6242 1588 6276
rect 122 6156 138 6190
rect 1572 6156 1588 6190
rect 122 6070 138 6104
rect 1572 6070 1588 6104
rect 122 5984 138 6018
rect 1572 5984 1588 6018
rect 122 5898 138 5932
rect 1572 5898 1588 5932
rect 122 5812 138 5846
rect 1572 5812 1588 5846
rect 122 5726 138 5760
rect 1572 5726 1588 5760
rect 122 5640 138 5674
rect 1572 5640 1588 5674
rect 122 5554 138 5588
rect 1572 5554 1588 5588
rect 122 5468 138 5502
rect 1572 5468 1588 5502
rect 122 5382 138 5416
rect 1572 5382 1588 5416
rect 122 5296 138 5330
rect 1572 5296 1588 5330
rect 122 5210 138 5244
rect 1572 5210 1588 5244
rect 122 5124 138 5158
rect 1572 5124 1588 5158
rect 122 5038 138 5072
rect 1572 5038 1588 5072
rect 122 4952 138 4986
rect 1572 4952 1588 4986
rect 122 4866 138 4900
rect 1572 4866 1588 4900
rect 122 4780 138 4814
rect 1572 4780 1588 4814
rect 122 4694 138 4728
rect 1572 4694 1588 4728
rect 122 4608 138 4642
rect 1572 4608 1588 4642
rect 122 4522 138 4556
rect 1572 4522 1588 4556
rect 122 4436 138 4470
rect 1572 4436 1588 4470
rect 122 4350 138 4384
rect 1572 4350 1588 4384
rect 122 4264 138 4298
rect 1572 4264 1588 4298
rect 122 4178 138 4212
rect 1572 4178 1588 4212
rect 122 4092 138 4126
rect 1572 4092 1588 4126
rect 122 4006 138 4040
rect 1572 4006 1588 4040
rect 122 3920 138 3954
rect 1572 3920 1588 3954
rect 122 3834 138 3868
rect 1572 3834 1588 3868
rect 122 3748 138 3782
rect 1572 3748 1588 3782
rect 122 3662 138 3696
rect 1572 3662 1588 3696
rect 122 3576 138 3610
rect 1572 3576 1588 3610
rect 122 3490 138 3524
rect 1572 3490 1588 3524
rect 122 3404 138 3438
rect 1572 3404 1588 3438
rect 122 3318 138 3352
rect 1572 3318 1588 3352
rect 122 3232 138 3266
rect 1572 3232 1588 3266
rect 122 3146 138 3180
rect 1572 3146 1588 3180
rect 122 3060 138 3094
rect 1572 3060 1588 3094
rect 122 2974 138 3008
rect 1572 2974 1588 3008
rect 122 2888 138 2922
rect 1572 2888 1588 2922
rect 122 2802 138 2836
rect 1572 2802 1588 2836
rect 122 2716 138 2750
rect 1572 2716 1588 2750
rect 122 2630 138 2664
rect 1572 2630 1588 2664
rect 122 2544 138 2578
rect 1572 2544 1588 2578
rect 122 2458 138 2492
rect 1572 2458 1588 2492
rect 122 2372 138 2406
rect 1572 2372 1588 2406
rect 122 2286 138 2320
rect 1572 2286 1588 2320
rect 122 2200 138 2234
rect 1572 2200 1588 2234
rect 122 2114 138 2148
rect 1572 2114 1588 2148
rect 122 2028 138 2062
rect 1572 2028 1588 2062
rect 122 1942 138 1976
rect 1572 1942 1588 1976
rect 122 1856 138 1890
rect 1572 1856 1588 1890
rect 122 1770 138 1804
rect 1572 1770 1588 1804
rect 122 1684 138 1718
rect 1572 1684 1588 1718
rect 122 1598 138 1632
rect 1572 1598 1588 1632
rect 122 1512 138 1546
rect 1572 1512 1588 1546
rect 122 1426 138 1460
rect 1572 1426 1588 1460
rect 122 1340 138 1374
rect 1572 1340 1588 1374
rect 122 1254 138 1288
rect 1572 1254 1588 1288
rect 122 1168 138 1202
rect 1572 1168 1588 1202
rect 122 1082 138 1116
rect 1572 1082 1588 1116
rect 122 996 138 1030
rect 1572 996 1588 1030
rect 122 910 138 944
rect 1572 910 1588 944
rect 122 824 138 858
rect 1572 824 1588 858
rect 122 738 138 772
rect 1572 738 1588 772
rect 122 652 138 686
rect 1572 652 1588 686
rect 122 566 138 600
rect 1572 566 1588 600
rect 122 480 138 514
rect 1572 480 1588 514
rect 122 394 138 428
rect 1572 394 1588 428
rect 122 308 138 342
rect 1572 308 1588 342
rect 122 222 138 256
rect 1572 222 1588 256
rect 122 136 138 170
rect 1572 136 1588 170
rect 1628 163 1662 179
rect 36 70 70 100
rect 1710 70 1744 100
rect 36 36 100 70
rect 1680 36 1744 70
<< viali >>
rect 100 21220 1680 21254
rect 36 100 70 21190
rect 138 21120 1572 21154
rect 138 21034 1572 21068
rect 138 20948 1572 20982
rect 138 20862 1572 20896
rect 138 20776 1572 20810
rect 138 20690 1572 20724
rect 138 20604 1572 20638
rect 138 20518 1572 20552
rect 138 20432 1572 20466
rect 138 20346 1572 20380
rect 138 20260 1572 20294
rect 138 20174 1572 20208
rect 138 20088 1572 20122
rect 138 20002 1572 20036
rect 138 19916 1572 19950
rect 138 19830 1572 19864
rect 138 19744 1572 19778
rect 138 19658 1572 19692
rect 138 19572 1572 19606
rect 138 19486 1572 19520
rect 138 19400 1572 19434
rect 138 19314 1572 19348
rect 138 19228 1572 19262
rect 138 19142 1572 19176
rect 138 19056 1572 19090
rect 138 18970 1572 19004
rect 138 18884 1572 18918
rect 138 18798 1572 18832
rect 138 18712 1572 18746
rect 138 18626 1572 18660
rect 138 18540 1572 18574
rect 138 18454 1572 18488
rect 138 18368 1572 18402
rect 138 18282 1572 18316
rect 138 18196 1572 18230
rect 138 18110 1572 18144
rect 138 18024 1572 18058
rect 138 17938 1572 17972
rect 138 17852 1572 17886
rect 138 17766 1572 17800
rect 138 17680 1572 17714
rect 138 17594 1572 17628
rect 138 17508 1572 17542
rect 138 17422 1572 17456
rect 138 17336 1572 17370
rect 138 17250 1572 17284
rect 138 17164 1572 17198
rect 138 17078 1572 17112
rect 138 16992 1572 17026
rect 138 16906 1572 16940
rect 138 16820 1572 16854
rect 138 16734 1572 16768
rect 138 16648 1572 16682
rect 138 16562 1572 16596
rect 138 16476 1572 16510
rect 138 16390 1572 16424
rect 138 16304 1572 16338
rect 138 16218 1572 16252
rect 138 16132 1572 16166
rect 138 16046 1572 16080
rect 138 15960 1572 15994
rect 138 15874 1572 15908
rect 138 15788 1572 15822
rect 138 15702 1572 15736
rect 138 15616 1572 15650
rect 138 15530 1572 15564
rect 138 15444 1572 15478
rect 138 15358 1572 15392
rect 138 15272 1572 15306
rect 138 15186 1572 15220
rect 138 15100 1572 15134
rect 138 15014 1572 15048
rect 138 14928 1572 14962
rect 138 14842 1572 14876
rect 138 14756 1572 14790
rect 138 14670 1572 14704
rect 138 14584 1572 14618
rect 138 14498 1572 14532
rect 138 14412 1572 14446
rect 138 14326 1572 14360
rect 138 14240 1572 14274
rect 138 14154 1572 14188
rect 138 14068 1572 14102
rect 138 13982 1572 14016
rect 138 13896 1572 13930
rect 138 13810 1572 13844
rect 138 13724 1572 13758
rect 138 13638 1572 13672
rect 138 13552 1572 13586
rect 138 13466 1572 13500
rect 138 13380 1572 13414
rect 138 13294 1572 13328
rect 138 13208 1572 13242
rect 138 13122 1572 13156
rect 138 13036 1572 13070
rect 138 12950 1572 12984
rect 138 12864 1572 12898
rect 138 12778 1572 12812
rect 138 12692 1572 12726
rect 138 12606 1572 12640
rect 138 12520 1572 12554
rect 138 12434 1572 12468
rect 138 12348 1572 12382
rect 138 12262 1572 12296
rect 138 12176 1572 12210
rect 138 12090 1572 12124
rect 138 12004 1572 12038
rect 138 11918 1572 11952
rect 138 11832 1572 11866
rect 138 11746 1572 11780
rect 138 11660 1572 11694
rect 138 11574 1572 11608
rect 138 11488 1572 11522
rect 138 11402 1572 11436
rect 138 11316 1572 11350
rect 138 11230 1572 11264
rect 138 11144 1572 11178
rect 138 11058 1572 11092
rect 138 10972 1572 11006
rect 138 10886 1572 10920
rect 138 10800 1572 10834
rect 138 10714 1572 10748
rect 138 10628 1572 10662
rect 138 10542 1572 10576
rect 138 10456 1572 10490
rect 138 10370 1572 10404
rect 138 10284 1572 10318
rect 138 10198 1572 10232
rect 138 10112 1572 10146
rect 138 10026 1572 10060
rect 138 9940 1572 9974
rect 138 9854 1572 9888
rect 138 9768 1572 9802
rect 138 9682 1572 9716
rect 138 9596 1572 9630
rect 138 9510 1572 9544
rect 138 9424 1572 9458
rect 138 9338 1572 9372
rect 138 9252 1572 9286
rect 138 9166 1572 9200
rect 138 9080 1572 9114
rect 138 8994 1572 9028
rect 138 8908 1572 8942
rect 138 8822 1572 8856
rect 138 8736 1572 8770
rect 138 8650 1572 8684
rect 138 8564 1572 8598
rect 138 8478 1572 8512
rect 138 8392 1572 8426
rect 138 8306 1572 8340
rect 138 8220 1572 8254
rect 138 8134 1572 8168
rect 138 8048 1572 8082
rect 138 7962 1572 7996
rect 138 7876 1572 7910
rect 138 7790 1572 7824
rect 138 7704 1572 7738
rect 138 7618 1572 7652
rect 138 7532 1572 7566
rect 138 7446 1572 7480
rect 138 7360 1572 7394
rect 138 7274 1572 7308
rect 138 7188 1572 7222
rect 138 7102 1572 7136
rect 138 7016 1572 7050
rect 138 6930 1572 6964
rect 138 6844 1572 6878
rect 138 6758 1572 6792
rect 138 6672 1572 6706
rect 138 6586 1572 6620
rect 138 6500 1572 6534
rect 138 6414 1572 6448
rect 138 6328 1572 6362
rect 138 6242 1572 6276
rect 138 6156 1572 6190
rect 138 6070 1572 6104
rect 138 5984 1572 6018
rect 138 5898 1572 5932
rect 138 5812 1572 5846
rect 138 5726 1572 5760
rect 138 5640 1572 5674
rect 138 5554 1572 5588
rect 138 5468 1572 5502
rect 138 5382 1572 5416
rect 138 5296 1572 5330
rect 138 5210 1572 5244
rect 138 5124 1572 5158
rect 138 5038 1572 5072
rect 138 4952 1572 4986
rect 138 4866 1572 4900
rect 138 4780 1572 4814
rect 138 4694 1572 4728
rect 138 4608 1572 4642
rect 138 4522 1572 4556
rect 138 4436 1572 4470
rect 138 4350 1572 4384
rect 138 4264 1572 4298
rect 138 4178 1572 4212
rect 138 4092 1572 4126
rect 138 4006 1572 4040
rect 138 3920 1572 3954
rect 138 3834 1572 3868
rect 138 3748 1572 3782
rect 138 3662 1572 3696
rect 138 3576 1572 3610
rect 138 3490 1572 3524
rect 138 3404 1572 3438
rect 138 3318 1572 3352
rect 138 3232 1572 3266
rect 138 3146 1572 3180
rect 138 3060 1572 3094
rect 138 2974 1572 3008
rect 138 2888 1572 2922
rect 138 2802 1572 2836
rect 138 2716 1572 2750
rect 138 2630 1572 2664
rect 138 2544 1572 2578
rect 138 2458 1572 2492
rect 138 2372 1572 2406
rect 138 2286 1572 2320
rect 138 2200 1572 2234
rect 138 2114 1572 2148
rect 138 2028 1572 2062
rect 138 1942 1572 1976
rect 138 1856 1572 1890
rect 138 1770 1572 1804
rect 138 1684 1572 1718
rect 138 1598 1572 1632
rect 138 1512 1572 1546
rect 138 1426 1572 1460
rect 138 1340 1572 1374
rect 138 1254 1572 1288
rect 138 1168 1572 1202
rect 138 1082 1572 1116
rect 138 996 1572 1030
rect 138 910 1572 944
rect 138 824 1572 858
rect 138 738 1572 772
rect 138 652 1572 686
rect 138 566 1572 600
rect 138 480 1572 514
rect 138 394 1572 428
rect 138 308 1572 342
rect 138 222 1572 256
rect 1628 179 1662 21111
rect 138 136 1572 170
rect 1710 100 1744 21190
rect 100 36 1680 70
<< metal1 >>
rect 30 21254 1750 21260
rect 30 21220 100 21254
rect 1680 21220 1750 21254
rect 30 21214 1750 21220
rect 30 21190 76 21214
rect 30 100 36 21190
rect 70 100 76 21190
rect 1704 21190 1750 21214
rect 894 21160 900 21163
rect 126 21154 900 21160
rect 1548 21160 1554 21163
rect 1548 21154 1584 21160
rect 126 21120 138 21154
rect 1572 21120 1584 21154
rect 126 21114 900 21120
rect 894 21111 900 21114
rect 1548 21114 1584 21120
rect 1618 21121 1672 21127
rect 1548 21111 1554 21114
rect 156 21074 162 21077
rect 126 21068 162 21074
rect 810 21074 816 21077
rect 810 21068 1584 21074
rect 126 21034 138 21068
rect 1572 21034 1584 21068
rect 126 21028 162 21034
rect 156 21025 162 21028
rect 810 21028 1584 21034
rect 810 21025 816 21028
rect 894 20988 900 20991
rect 126 20982 900 20988
rect 1548 20988 1554 20991
rect 1548 20982 1584 20988
rect 126 20948 138 20982
rect 1572 20948 1584 20982
rect 126 20942 900 20948
rect 894 20939 900 20942
rect 1548 20942 1584 20948
rect 1548 20939 1554 20942
rect 156 20902 162 20905
rect 126 20896 162 20902
rect 810 20902 816 20905
rect 810 20896 1584 20902
rect 126 20862 138 20896
rect 1572 20862 1584 20896
rect 126 20856 162 20862
rect 156 20853 162 20856
rect 810 20856 1584 20862
rect 810 20853 816 20856
rect 894 20816 900 20819
rect 126 20810 900 20816
rect 1548 20816 1554 20819
rect 1548 20810 1584 20816
rect 126 20776 138 20810
rect 1572 20776 1584 20810
rect 126 20770 900 20776
rect 894 20767 900 20770
rect 1548 20770 1584 20776
rect 1548 20767 1554 20770
rect 156 20730 162 20733
rect 126 20724 162 20730
rect 810 20730 816 20733
rect 810 20724 1584 20730
rect 126 20690 138 20724
rect 1572 20690 1584 20724
rect 126 20684 162 20690
rect 156 20681 162 20684
rect 810 20684 1584 20690
rect 810 20681 816 20684
rect 894 20644 900 20647
rect 126 20638 900 20644
rect 1548 20644 1554 20647
rect 1548 20638 1584 20644
rect 126 20604 138 20638
rect 1572 20604 1584 20638
rect 126 20598 900 20604
rect 894 20595 900 20598
rect 1548 20598 1584 20604
rect 1548 20595 1554 20598
rect 156 20558 162 20561
rect 126 20552 162 20558
rect 810 20558 816 20561
rect 810 20552 1584 20558
rect 126 20518 138 20552
rect 1572 20518 1584 20552
rect 126 20512 162 20518
rect 156 20509 162 20512
rect 810 20512 1584 20518
rect 810 20509 816 20512
rect 894 20472 900 20475
rect 126 20466 900 20472
rect 1548 20472 1554 20475
rect 1548 20466 1584 20472
rect 126 20432 138 20466
rect 1572 20432 1584 20466
rect 126 20426 900 20432
rect 894 20423 900 20426
rect 1548 20426 1584 20432
rect 1548 20423 1554 20426
rect 156 20386 162 20389
rect 126 20380 162 20386
rect 810 20386 816 20389
rect 810 20380 1584 20386
rect 126 20346 138 20380
rect 1572 20346 1584 20380
rect 126 20340 162 20346
rect 156 20337 162 20340
rect 810 20340 1584 20346
rect 810 20337 816 20340
rect 894 20300 900 20303
rect 126 20294 900 20300
rect 1548 20300 1554 20303
rect 1548 20294 1584 20300
rect 126 20260 138 20294
rect 1572 20260 1584 20294
rect 126 20254 900 20260
rect 894 20251 900 20254
rect 1548 20254 1584 20260
rect 1548 20251 1554 20254
rect 156 20214 162 20217
rect 126 20208 162 20214
rect 810 20214 816 20217
rect 810 20208 1584 20214
rect 126 20174 138 20208
rect 1572 20174 1584 20208
rect 126 20168 162 20174
rect 156 20165 162 20168
rect 810 20168 1584 20174
rect 810 20165 816 20168
rect 894 20128 900 20131
rect 126 20122 900 20128
rect 1548 20128 1554 20131
rect 1548 20122 1584 20128
rect 126 20088 138 20122
rect 1572 20088 1584 20122
rect 126 20082 900 20088
rect 894 20079 900 20082
rect 1548 20082 1584 20088
rect 1548 20079 1554 20082
rect 156 20042 162 20045
rect 126 20036 162 20042
rect 810 20042 816 20045
rect 810 20036 1584 20042
rect 126 20002 138 20036
rect 1572 20002 1584 20036
rect 126 19996 162 20002
rect 156 19993 162 19996
rect 810 19996 1584 20002
rect 810 19993 816 19996
rect 894 19956 900 19959
rect 126 19950 900 19956
rect 1548 19956 1554 19959
rect 1548 19950 1584 19956
rect 126 19916 138 19950
rect 1572 19916 1584 19950
rect 126 19910 900 19916
rect 894 19907 900 19910
rect 1548 19910 1584 19916
rect 1548 19907 1554 19910
rect 156 19870 162 19873
rect 126 19864 162 19870
rect 810 19870 816 19873
rect 810 19864 1584 19870
rect 126 19830 138 19864
rect 1572 19830 1584 19864
rect 126 19824 162 19830
rect 156 19821 162 19824
rect 810 19824 1584 19830
rect 810 19821 816 19824
rect 894 19784 900 19787
rect 126 19778 900 19784
rect 1548 19784 1554 19787
rect 1548 19778 1584 19784
rect 126 19744 138 19778
rect 1572 19744 1584 19778
rect 126 19738 900 19744
rect 894 19735 900 19738
rect 1548 19738 1584 19744
rect 1548 19735 1554 19738
rect 156 19698 162 19701
rect 126 19692 162 19698
rect 810 19698 816 19701
rect 810 19692 1584 19698
rect 126 19658 138 19692
rect 1572 19658 1584 19692
rect 126 19652 162 19658
rect 156 19649 162 19652
rect 810 19652 1584 19658
rect 810 19649 816 19652
rect 894 19612 900 19615
rect 126 19606 900 19612
rect 1548 19612 1554 19615
rect 1548 19606 1584 19612
rect 126 19572 138 19606
rect 1572 19572 1584 19606
rect 126 19566 900 19572
rect 894 19563 900 19566
rect 1548 19566 1584 19572
rect 1548 19563 1554 19566
rect 156 19526 162 19529
rect 126 19520 162 19526
rect 810 19526 816 19529
rect 810 19520 1584 19526
rect 126 19486 138 19520
rect 1572 19486 1584 19520
rect 126 19480 162 19486
rect 156 19477 162 19480
rect 810 19480 1584 19486
rect 810 19477 816 19480
rect 894 19440 900 19443
rect 126 19434 900 19440
rect 1548 19440 1554 19443
rect 1548 19434 1584 19440
rect 126 19400 138 19434
rect 1572 19400 1584 19434
rect 126 19394 900 19400
rect 894 19391 900 19394
rect 1548 19394 1584 19400
rect 1548 19391 1554 19394
rect 156 19354 162 19357
rect 126 19348 162 19354
rect 810 19354 816 19357
rect 810 19348 1584 19354
rect 126 19314 138 19348
rect 1572 19314 1584 19348
rect 126 19308 162 19314
rect 156 19305 162 19308
rect 810 19308 1584 19314
rect 810 19305 816 19308
rect 894 19268 900 19271
rect 126 19262 900 19268
rect 1548 19268 1554 19271
rect 1548 19262 1584 19268
rect 126 19228 138 19262
rect 1572 19228 1584 19262
rect 126 19222 900 19228
rect 894 19219 900 19222
rect 1548 19222 1584 19228
rect 1548 19219 1554 19222
rect 156 19182 162 19185
rect 126 19176 162 19182
rect 810 19182 816 19185
rect 810 19176 1584 19182
rect 126 19142 138 19176
rect 1572 19142 1584 19176
rect 126 19136 162 19142
rect 156 19133 162 19136
rect 810 19136 1584 19142
rect 810 19133 816 19136
rect 894 19096 900 19099
rect 126 19090 900 19096
rect 1548 19096 1554 19099
rect 1548 19090 1584 19096
rect 126 19056 138 19090
rect 1572 19056 1584 19090
rect 126 19050 900 19056
rect 894 19047 900 19050
rect 1548 19050 1584 19056
rect 1548 19047 1554 19050
rect 156 19010 162 19013
rect 126 19004 162 19010
rect 810 19010 816 19013
rect 810 19004 1584 19010
rect 126 18970 138 19004
rect 1572 18970 1584 19004
rect 126 18964 162 18970
rect 156 18961 162 18964
rect 810 18964 1584 18970
rect 810 18961 816 18964
rect 894 18924 900 18927
rect 126 18918 900 18924
rect 1548 18924 1554 18927
rect 1548 18918 1584 18924
rect 126 18884 138 18918
rect 1572 18884 1584 18918
rect 126 18878 900 18884
rect 894 18875 900 18878
rect 1548 18878 1584 18884
rect 1548 18875 1554 18878
rect 156 18838 162 18841
rect 126 18832 162 18838
rect 810 18838 816 18841
rect 810 18832 1584 18838
rect 126 18798 138 18832
rect 1572 18798 1584 18832
rect 126 18792 162 18798
rect 156 18789 162 18792
rect 810 18792 1584 18798
rect 810 18789 816 18792
rect 894 18752 900 18755
rect 126 18746 900 18752
rect 1548 18752 1554 18755
rect 1548 18746 1584 18752
rect 126 18712 138 18746
rect 1572 18712 1584 18746
rect 126 18706 900 18712
rect 894 18703 900 18706
rect 1548 18706 1584 18712
rect 1548 18703 1554 18706
rect 156 18666 162 18669
rect 126 18660 162 18666
rect 810 18666 816 18669
rect 810 18660 1584 18666
rect 126 18626 138 18660
rect 1572 18626 1584 18660
rect 126 18620 162 18626
rect 156 18617 162 18620
rect 810 18620 1584 18626
rect 810 18617 816 18620
rect 894 18580 900 18583
rect 126 18574 900 18580
rect 1548 18580 1554 18583
rect 1548 18574 1584 18580
rect 126 18540 138 18574
rect 1572 18540 1584 18574
rect 126 18534 900 18540
rect 894 18531 900 18534
rect 1548 18534 1584 18540
rect 1548 18531 1554 18534
rect 156 18494 162 18497
rect 126 18488 162 18494
rect 810 18494 816 18497
rect 810 18488 1584 18494
rect 126 18454 138 18488
rect 1572 18454 1584 18488
rect 126 18448 162 18454
rect 156 18445 162 18448
rect 810 18448 1584 18454
rect 810 18445 816 18448
rect 894 18408 900 18411
rect 126 18402 900 18408
rect 1548 18408 1554 18411
rect 1548 18402 1584 18408
rect 126 18368 138 18402
rect 1572 18368 1584 18402
rect 126 18362 900 18368
rect 894 18359 900 18362
rect 1548 18362 1584 18368
rect 1548 18359 1554 18362
rect 156 18322 162 18325
rect 126 18316 162 18322
rect 810 18322 816 18325
rect 810 18316 1584 18322
rect 126 18282 138 18316
rect 1572 18282 1584 18316
rect 126 18276 162 18282
rect 156 18273 162 18276
rect 810 18276 1584 18282
rect 810 18273 816 18276
rect 894 18236 900 18239
rect 126 18230 900 18236
rect 1548 18236 1554 18239
rect 1548 18230 1584 18236
rect 126 18196 138 18230
rect 1572 18196 1584 18230
rect 126 18190 900 18196
rect 894 18187 900 18190
rect 1548 18190 1584 18196
rect 1548 18187 1554 18190
rect 156 18150 162 18153
rect 126 18144 162 18150
rect 810 18150 816 18153
rect 810 18144 1584 18150
rect 126 18110 138 18144
rect 1572 18110 1584 18144
rect 126 18104 162 18110
rect 156 18101 162 18104
rect 810 18104 1584 18110
rect 810 18101 816 18104
rect 894 18064 900 18067
rect 126 18058 900 18064
rect 1548 18064 1554 18067
rect 1548 18058 1584 18064
rect 126 18024 138 18058
rect 1572 18024 1584 18058
rect 126 18018 900 18024
rect 894 18015 900 18018
rect 1548 18018 1584 18024
rect 1548 18015 1554 18018
rect 156 17978 162 17981
rect 126 17972 162 17978
rect 810 17978 816 17981
rect 810 17972 1584 17978
rect 126 17938 138 17972
rect 1572 17938 1584 17972
rect 126 17932 162 17938
rect 156 17929 162 17932
rect 810 17932 1584 17938
rect 810 17929 816 17932
rect 894 17892 900 17895
rect 126 17886 900 17892
rect 1548 17892 1554 17895
rect 1548 17886 1584 17892
rect 126 17852 138 17886
rect 1572 17852 1584 17886
rect 126 17846 900 17852
rect 894 17843 900 17846
rect 1548 17846 1584 17852
rect 1548 17843 1554 17846
rect 156 17806 162 17809
rect 126 17800 162 17806
rect 810 17806 816 17809
rect 810 17800 1584 17806
rect 126 17766 138 17800
rect 1572 17766 1584 17800
rect 126 17760 162 17766
rect 156 17757 162 17760
rect 810 17760 1584 17766
rect 810 17757 816 17760
rect 894 17720 900 17723
rect 126 17714 900 17720
rect 1548 17720 1554 17723
rect 1548 17714 1584 17720
rect 126 17680 138 17714
rect 1572 17680 1584 17714
rect 126 17674 900 17680
rect 894 17671 900 17674
rect 1548 17674 1584 17680
rect 1548 17671 1554 17674
rect 156 17634 162 17637
rect 126 17628 162 17634
rect 810 17634 816 17637
rect 810 17628 1584 17634
rect 126 17594 138 17628
rect 1572 17594 1584 17628
rect 126 17588 162 17594
rect 156 17585 162 17588
rect 810 17588 1584 17594
rect 810 17585 816 17588
rect 894 17548 900 17551
rect 126 17542 900 17548
rect 1548 17548 1554 17551
rect 1548 17542 1584 17548
rect 126 17508 138 17542
rect 1572 17508 1584 17542
rect 126 17502 900 17508
rect 894 17499 900 17502
rect 1548 17502 1584 17508
rect 1548 17499 1554 17502
rect 156 17462 162 17465
rect 126 17456 162 17462
rect 810 17462 816 17465
rect 810 17456 1584 17462
rect 126 17422 138 17456
rect 1572 17422 1584 17456
rect 126 17416 162 17422
rect 156 17413 162 17416
rect 810 17416 1584 17422
rect 810 17413 816 17416
rect 894 17376 900 17379
rect 126 17370 900 17376
rect 1548 17376 1554 17379
rect 1548 17370 1584 17376
rect 126 17336 138 17370
rect 1572 17336 1584 17370
rect 126 17330 900 17336
rect 894 17327 900 17330
rect 1548 17330 1584 17336
rect 1548 17327 1554 17330
rect 156 17290 162 17293
rect 126 17284 162 17290
rect 810 17290 816 17293
rect 810 17284 1584 17290
rect 126 17250 138 17284
rect 1572 17250 1584 17284
rect 126 17244 162 17250
rect 156 17241 162 17244
rect 810 17244 1584 17250
rect 810 17241 816 17244
rect 894 17204 900 17207
rect 126 17198 900 17204
rect 1548 17204 1554 17207
rect 1548 17198 1584 17204
rect 126 17164 138 17198
rect 1572 17164 1584 17198
rect 126 17158 900 17164
rect 894 17155 900 17158
rect 1548 17158 1584 17164
rect 1548 17155 1554 17158
rect 156 17118 162 17121
rect 126 17112 162 17118
rect 810 17118 816 17121
rect 810 17112 1584 17118
rect 126 17078 138 17112
rect 1572 17078 1584 17112
rect 126 17072 162 17078
rect 156 17069 162 17072
rect 810 17072 1584 17078
rect 810 17069 816 17072
rect 894 17032 900 17035
rect 126 17026 900 17032
rect 1548 17032 1554 17035
rect 1548 17026 1584 17032
rect 126 16992 138 17026
rect 1572 16992 1584 17026
rect 126 16986 900 16992
rect 894 16983 900 16986
rect 1548 16986 1584 16992
rect 1548 16983 1554 16986
rect 156 16946 162 16949
rect 126 16940 162 16946
rect 810 16946 816 16949
rect 810 16940 1584 16946
rect 126 16906 138 16940
rect 1572 16906 1584 16940
rect 126 16900 162 16906
rect 156 16897 162 16900
rect 810 16900 1584 16906
rect 810 16897 816 16900
rect 894 16860 900 16863
rect 126 16854 900 16860
rect 1548 16860 1554 16863
rect 1548 16854 1584 16860
rect 126 16820 138 16854
rect 1572 16820 1584 16854
rect 126 16814 900 16820
rect 894 16811 900 16814
rect 1548 16814 1584 16820
rect 1548 16811 1554 16814
rect 156 16774 162 16777
rect 126 16768 162 16774
rect 810 16774 816 16777
rect 810 16768 1584 16774
rect 126 16734 138 16768
rect 1572 16734 1584 16768
rect 126 16728 162 16734
rect 156 16725 162 16728
rect 810 16728 1584 16734
rect 810 16725 816 16728
rect 894 16688 900 16691
rect 126 16682 900 16688
rect 1548 16688 1554 16691
rect 1548 16682 1584 16688
rect 126 16648 138 16682
rect 1572 16648 1584 16682
rect 126 16642 900 16648
rect 894 16639 900 16642
rect 1548 16642 1584 16648
rect 1548 16639 1554 16642
rect 156 16602 162 16605
rect 126 16596 162 16602
rect 810 16602 816 16605
rect 810 16596 1584 16602
rect 126 16562 138 16596
rect 1572 16562 1584 16596
rect 126 16556 162 16562
rect 156 16553 162 16556
rect 810 16556 1584 16562
rect 810 16553 816 16556
rect 894 16516 900 16519
rect 126 16510 900 16516
rect 1548 16516 1554 16519
rect 1548 16510 1584 16516
rect 126 16476 138 16510
rect 1572 16476 1584 16510
rect 126 16470 900 16476
rect 894 16467 900 16470
rect 1548 16470 1584 16476
rect 1548 16467 1554 16470
rect 156 16430 162 16433
rect 126 16424 162 16430
rect 810 16430 816 16433
rect 810 16424 1584 16430
rect 126 16390 138 16424
rect 1572 16390 1584 16424
rect 126 16384 162 16390
rect 156 16381 162 16384
rect 810 16384 1584 16390
rect 810 16381 816 16384
rect 894 16344 900 16347
rect 126 16338 900 16344
rect 1548 16344 1554 16347
rect 1548 16338 1584 16344
rect 126 16304 138 16338
rect 1572 16304 1584 16338
rect 126 16298 900 16304
rect 894 16295 900 16298
rect 1548 16298 1584 16304
rect 1548 16295 1554 16298
rect 156 16258 162 16261
rect 126 16252 162 16258
rect 810 16258 816 16261
rect 810 16252 1584 16258
rect 126 16218 138 16252
rect 1572 16218 1584 16252
rect 126 16212 162 16218
rect 156 16209 162 16212
rect 810 16212 1584 16218
rect 810 16209 816 16212
rect 894 16172 900 16175
rect 126 16166 900 16172
rect 1548 16172 1554 16175
rect 1548 16166 1584 16172
rect 126 16132 138 16166
rect 1572 16132 1584 16166
rect 126 16126 900 16132
rect 894 16123 900 16126
rect 1548 16126 1584 16132
rect 1548 16123 1554 16126
rect 156 16086 162 16089
rect 126 16080 162 16086
rect 810 16086 816 16089
rect 810 16080 1584 16086
rect 126 16046 138 16080
rect 1572 16046 1584 16080
rect 126 16040 162 16046
rect 156 16037 162 16040
rect 810 16040 1584 16046
rect 810 16037 816 16040
rect 894 16000 900 16003
rect 126 15994 900 16000
rect 1548 16000 1554 16003
rect 1548 15994 1584 16000
rect 126 15960 138 15994
rect 1572 15960 1584 15994
rect 126 15954 900 15960
rect 894 15951 900 15954
rect 1548 15954 1584 15960
rect 1548 15951 1554 15954
rect 156 15914 162 15917
rect 126 15908 162 15914
rect 810 15914 816 15917
rect 810 15908 1584 15914
rect 126 15874 138 15908
rect 1572 15874 1584 15908
rect 126 15868 162 15874
rect 156 15865 162 15868
rect 810 15868 1584 15874
rect 810 15865 816 15868
rect 894 15828 900 15831
rect 126 15822 900 15828
rect 1548 15828 1554 15831
rect 1548 15822 1584 15828
rect 126 15788 138 15822
rect 1572 15788 1584 15822
rect 126 15782 900 15788
rect 894 15779 900 15782
rect 1548 15782 1584 15788
rect 1548 15779 1554 15782
rect 156 15742 162 15745
rect 126 15736 162 15742
rect 810 15742 816 15745
rect 810 15736 1584 15742
rect 126 15702 138 15736
rect 1572 15702 1584 15736
rect 126 15696 162 15702
rect 156 15693 162 15696
rect 810 15696 1584 15702
rect 810 15693 816 15696
rect 894 15656 900 15659
rect 126 15650 900 15656
rect 1548 15656 1554 15659
rect 1548 15650 1584 15656
rect 126 15616 138 15650
rect 1572 15616 1584 15650
rect 126 15610 900 15616
rect 894 15607 900 15610
rect 1548 15610 1584 15616
rect 1548 15607 1554 15610
rect 156 15570 162 15573
rect 126 15564 162 15570
rect 810 15570 816 15573
rect 810 15564 1584 15570
rect 126 15530 138 15564
rect 1572 15530 1584 15564
rect 126 15524 162 15530
rect 156 15521 162 15524
rect 810 15524 1584 15530
rect 810 15521 816 15524
rect 894 15484 900 15487
rect 126 15478 900 15484
rect 1548 15484 1554 15487
rect 1548 15478 1584 15484
rect 126 15444 138 15478
rect 1572 15444 1584 15478
rect 126 15438 900 15444
rect 894 15435 900 15438
rect 1548 15438 1584 15444
rect 1548 15435 1554 15438
rect 156 15398 162 15401
rect 126 15392 162 15398
rect 810 15398 816 15401
rect 810 15392 1584 15398
rect 126 15358 138 15392
rect 1572 15358 1584 15392
rect 126 15352 162 15358
rect 156 15349 162 15352
rect 810 15352 1584 15358
rect 810 15349 816 15352
rect 894 15312 900 15315
rect 126 15306 900 15312
rect 1548 15312 1554 15315
rect 1548 15306 1584 15312
rect 126 15272 138 15306
rect 1572 15272 1584 15306
rect 126 15266 900 15272
rect 894 15263 900 15266
rect 1548 15266 1584 15272
rect 1548 15263 1554 15266
rect 156 15226 162 15229
rect 126 15220 162 15226
rect 810 15226 816 15229
rect 810 15220 1584 15226
rect 126 15186 138 15220
rect 1572 15186 1584 15220
rect 126 15180 162 15186
rect 156 15177 162 15180
rect 810 15180 1584 15186
rect 810 15177 816 15180
rect 894 15140 900 15143
rect 126 15134 900 15140
rect 1548 15140 1554 15143
rect 1548 15134 1584 15140
rect 126 15100 138 15134
rect 1572 15100 1584 15134
rect 126 15094 900 15100
rect 894 15091 900 15094
rect 1548 15094 1584 15100
rect 1548 15091 1554 15094
rect 156 15054 162 15057
rect 126 15048 162 15054
rect 810 15054 816 15057
rect 810 15048 1584 15054
rect 126 15014 138 15048
rect 1572 15014 1584 15048
rect 126 15008 162 15014
rect 156 15005 162 15008
rect 810 15008 1584 15014
rect 810 15005 816 15008
rect 894 14968 900 14971
rect 126 14962 900 14968
rect 1548 14968 1554 14971
rect 1548 14962 1584 14968
rect 126 14928 138 14962
rect 1572 14928 1584 14962
rect 126 14922 900 14928
rect 894 14919 900 14922
rect 1548 14922 1584 14928
rect 1548 14919 1554 14922
rect 156 14882 162 14885
rect 126 14876 162 14882
rect 810 14882 816 14885
rect 810 14876 1584 14882
rect 126 14842 138 14876
rect 1572 14842 1584 14876
rect 126 14836 162 14842
rect 156 14833 162 14836
rect 810 14836 1584 14842
rect 810 14833 816 14836
rect 894 14796 900 14799
rect 126 14790 900 14796
rect 1548 14796 1554 14799
rect 1548 14790 1584 14796
rect 126 14756 138 14790
rect 1572 14756 1584 14790
rect 126 14750 900 14756
rect 894 14747 900 14750
rect 1548 14750 1584 14756
rect 1548 14747 1554 14750
rect 156 14710 162 14713
rect 126 14704 162 14710
rect 810 14710 816 14713
rect 810 14704 1584 14710
rect 126 14670 138 14704
rect 1572 14670 1584 14704
rect 126 14664 162 14670
rect 156 14661 162 14664
rect 810 14664 1584 14670
rect 810 14661 816 14664
rect 894 14624 900 14627
rect 126 14618 900 14624
rect 1548 14624 1554 14627
rect 1548 14618 1584 14624
rect 126 14584 138 14618
rect 1572 14584 1584 14618
rect 126 14578 900 14584
rect 894 14575 900 14578
rect 1548 14578 1584 14584
rect 1548 14575 1554 14578
rect 156 14538 162 14541
rect 126 14532 162 14538
rect 810 14538 816 14541
rect 810 14532 1584 14538
rect 126 14498 138 14532
rect 1572 14498 1584 14532
rect 126 14492 162 14498
rect 156 14489 162 14492
rect 810 14492 1584 14498
rect 810 14489 816 14492
rect 894 14452 900 14455
rect 126 14446 900 14452
rect 1548 14452 1554 14455
rect 1548 14446 1584 14452
rect 126 14412 138 14446
rect 1572 14412 1584 14446
rect 126 14406 900 14412
rect 894 14403 900 14406
rect 1548 14406 1584 14412
rect 1548 14403 1554 14406
rect 156 14366 162 14369
rect 126 14360 162 14366
rect 810 14366 816 14369
rect 810 14360 1584 14366
rect 126 14326 138 14360
rect 1572 14326 1584 14360
rect 126 14320 162 14326
rect 156 14317 162 14320
rect 810 14320 1584 14326
rect 810 14317 816 14320
rect 894 14280 900 14283
rect 126 14274 900 14280
rect 1548 14280 1554 14283
rect 1548 14274 1584 14280
rect 126 14240 138 14274
rect 1572 14240 1584 14274
rect 126 14234 900 14240
rect 894 14231 900 14234
rect 1548 14234 1584 14240
rect 1548 14231 1554 14234
rect 156 14194 162 14197
rect 126 14188 162 14194
rect 810 14194 816 14197
rect 810 14188 1584 14194
rect 126 14154 138 14188
rect 1572 14154 1584 14188
rect 126 14148 162 14154
rect 156 14145 162 14148
rect 810 14148 1584 14154
rect 810 14145 816 14148
rect 894 14108 900 14111
rect 126 14102 900 14108
rect 1548 14108 1554 14111
rect 1548 14102 1584 14108
rect 126 14068 138 14102
rect 1572 14068 1584 14102
rect 126 14062 900 14068
rect 894 14059 900 14062
rect 1548 14062 1584 14068
rect 1548 14059 1554 14062
rect 156 14022 162 14025
rect 126 14016 162 14022
rect 810 14022 816 14025
rect 810 14016 1584 14022
rect 126 13982 138 14016
rect 1572 13982 1584 14016
rect 126 13976 162 13982
rect 156 13973 162 13976
rect 810 13976 1584 13982
rect 810 13973 816 13976
rect 894 13936 900 13939
rect 126 13930 900 13936
rect 1548 13936 1554 13939
rect 1548 13930 1584 13936
rect 126 13896 138 13930
rect 1572 13896 1584 13930
rect 126 13890 900 13896
rect 894 13887 900 13890
rect 1548 13890 1584 13896
rect 1548 13887 1554 13890
rect 156 13850 162 13853
rect 126 13844 162 13850
rect 810 13850 816 13853
rect 810 13844 1584 13850
rect 126 13810 138 13844
rect 1572 13810 1584 13844
rect 126 13804 162 13810
rect 156 13801 162 13804
rect 810 13804 1584 13810
rect 810 13801 816 13804
rect 894 13764 900 13767
rect 126 13758 900 13764
rect 1548 13764 1554 13767
rect 1548 13758 1584 13764
rect 126 13724 138 13758
rect 1572 13724 1584 13758
rect 126 13718 900 13724
rect 894 13715 900 13718
rect 1548 13718 1584 13724
rect 1548 13715 1554 13718
rect 156 13678 162 13681
rect 126 13672 162 13678
rect 810 13678 816 13681
rect 810 13672 1584 13678
rect 126 13638 138 13672
rect 1572 13638 1584 13672
rect 126 13632 162 13638
rect 156 13629 162 13632
rect 810 13632 1584 13638
rect 810 13629 816 13632
rect 894 13592 900 13595
rect 126 13586 900 13592
rect 1548 13592 1554 13595
rect 1548 13586 1584 13592
rect 126 13552 138 13586
rect 1572 13552 1584 13586
rect 126 13546 900 13552
rect 894 13543 900 13546
rect 1548 13546 1584 13552
rect 1548 13543 1554 13546
rect 156 13506 162 13509
rect 126 13500 162 13506
rect 810 13506 816 13509
rect 810 13500 1584 13506
rect 126 13466 138 13500
rect 1572 13466 1584 13500
rect 126 13460 162 13466
rect 156 13457 162 13460
rect 810 13460 1584 13466
rect 810 13457 816 13460
rect 894 13420 900 13423
rect 126 13414 900 13420
rect 1548 13420 1554 13423
rect 1548 13414 1584 13420
rect 126 13380 138 13414
rect 1572 13380 1584 13414
rect 126 13374 900 13380
rect 894 13371 900 13374
rect 1548 13374 1584 13380
rect 1548 13371 1554 13374
rect 156 13334 162 13337
rect 126 13328 162 13334
rect 810 13334 816 13337
rect 810 13328 1584 13334
rect 126 13294 138 13328
rect 1572 13294 1584 13328
rect 126 13288 162 13294
rect 156 13285 162 13288
rect 810 13288 1584 13294
rect 810 13285 816 13288
rect 894 13248 900 13251
rect 126 13242 900 13248
rect 1548 13248 1554 13251
rect 1548 13242 1584 13248
rect 126 13208 138 13242
rect 1572 13208 1584 13242
rect 126 13202 900 13208
rect 894 13199 900 13202
rect 1548 13202 1584 13208
rect 1548 13199 1554 13202
rect 156 13162 162 13165
rect 126 13156 162 13162
rect 810 13162 816 13165
rect 810 13156 1584 13162
rect 126 13122 138 13156
rect 1572 13122 1584 13156
rect 126 13116 162 13122
rect 156 13113 162 13116
rect 810 13116 1584 13122
rect 810 13113 816 13116
rect 894 13076 900 13079
rect 126 13070 900 13076
rect 1548 13076 1554 13079
rect 1548 13070 1584 13076
rect 126 13036 138 13070
rect 1572 13036 1584 13070
rect 126 13030 900 13036
rect 894 13027 900 13030
rect 1548 13030 1584 13036
rect 1548 13027 1554 13030
rect 156 12990 162 12993
rect 126 12984 162 12990
rect 810 12990 816 12993
rect 810 12984 1584 12990
rect 126 12950 138 12984
rect 1572 12950 1584 12984
rect 126 12944 162 12950
rect 156 12941 162 12944
rect 810 12944 1584 12950
rect 810 12941 816 12944
rect 894 12904 900 12907
rect 126 12898 900 12904
rect 1548 12904 1554 12907
rect 1548 12898 1584 12904
rect 126 12864 138 12898
rect 1572 12864 1584 12898
rect 126 12858 900 12864
rect 894 12855 900 12858
rect 1548 12858 1584 12864
rect 1548 12855 1554 12858
rect 156 12818 162 12821
rect 126 12812 162 12818
rect 810 12818 816 12821
rect 810 12812 1584 12818
rect 126 12778 138 12812
rect 1572 12778 1584 12812
rect 126 12772 162 12778
rect 156 12769 162 12772
rect 810 12772 1584 12778
rect 810 12769 816 12772
rect 894 12732 900 12735
rect 126 12726 900 12732
rect 1548 12732 1554 12735
rect 1548 12726 1584 12732
rect 126 12692 138 12726
rect 1572 12692 1584 12726
rect 126 12686 900 12692
rect 894 12683 900 12686
rect 1548 12686 1584 12692
rect 1548 12683 1554 12686
rect 156 12646 162 12649
rect 126 12640 162 12646
rect 810 12646 816 12649
rect 810 12640 1584 12646
rect 126 12606 138 12640
rect 1572 12606 1584 12640
rect 126 12600 162 12606
rect 156 12597 162 12600
rect 810 12600 1584 12606
rect 810 12597 816 12600
rect 894 12560 900 12563
rect 126 12554 900 12560
rect 1548 12560 1554 12563
rect 1548 12554 1584 12560
rect 126 12520 138 12554
rect 1572 12520 1584 12554
rect 126 12514 900 12520
rect 894 12511 900 12514
rect 1548 12514 1584 12520
rect 1548 12511 1554 12514
rect 156 12474 162 12477
rect 126 12468 162 12474
rect 810 12474 816 12477
rect 810 12468 1584 12474
rect 126 12434 138 12468
rect 1572 12434 1584 12468
rect 126 12428 162 12434
rect 156 12425 162 12428
rect 810 12428 1584 12434
rect 810 12425 816 12428
rect 894 12388 900 12391
rect 126 12382 900 12388
rect 1548 12388 1554 12391
rect 1548 12382 1584 12388
rect 126 12348 138 12382
rect 1572 12348 1584 12382
rect 126 12342 900 12348
rect 894 12339 900 12342
rect 1548 12342 1584 12348
rect 1548 12339 1554 12342
rect 156 12302 162 12305
rect 126 12296 162 12302
rect 810 12302 816 12305
rect 810 12296 1584 12302
rect 126 12262 138 12296
rect 1572 12262 1584 12296
rect 126 12256 162 12262
rect 156 12253 162 12256
rect 810 12256 1584 12262
rect 810 12253 816 12256
rect 894 12216 900 12219
rect 126 12210 900 12216
rect 1548 12216 1554 12219
rect 1548 12210 1584 12216
rect 126 12176 138 12210
rect 1572 12176 1584 12210
rect 126 12170 900 12176
rect 894 12167 900 12170
rect 1548 12170 1584 12176
rect 1548 12167 1554 12170
rect 156 12130 162 12133
rect 126 12124 162 12130
rect 810 12130 816 12133
rect 810 12124 1584 12130
rect 126 12090 138 12124
rect 1572 12090 1584 12124
rect 126 12084 162 12090
rect 156 12081 162 12084
rect 810 12084 1584 12090
rect 810 12081 816 12084
rect 894 12044 900 12047
rect 126 12038 900 12044
rect 1548 12044 1554 12047
rect 1548 12038 1584 12044
rect 126 12004 138 12038
rect 1572 12004 1584 12038
rect 126 11998 900 12004
rect 894 11995 900 11998
rect 1548 11998 1584 12004
rect 1548 11995 1554 11998
rect 156 11958 162 11961
rect 126 11952 162 11958
rect 810 11958 816 11961
rect 810 11952 1584 11958
rect 126 11918 138 11952
rect 1572 11918 1584 11952
rect 126 11912 162 11918
rect 156 11909 162 11912
rect 810 11912 1584 11918
rect 810 11909 816 11912
rect 894 11872 900 11875
rect 126 11866 900 11872
rect 1548 11872 1554 11875
rect 1548 11866 1584 11872
rect 126 11832 138 11866
rect 1572 11832 1584 11866
rect 126 11826 900 11832
rect 894 11823 900 11826
rect 1548 11826 1584 11832
rect 1548 11823 1554 11826
rect 156 11786 162 11789
rect 126 11780 162 11786
rect 810 11786 816 11789
rect 810 11780 1584 11786
rect 126 11746 138 11780
rect 1572 11746 1584 11780
rect 126 11740 162 11746
rect 156 11737 162 11740
rect 810 11740 1584 11746
rect 810 11737 816 11740
rect 894 11700 900 11703
rect 126 11694 900 11700
rect 1548 11700 1554 11703
rect 1548 11694 1584 11700
rect 126 11660 138 11694
rect 1572 11660 1584 11694
rect 126 11654 900 11660
rect 894 11651 900 11654
rect 1548 11654 1584 11660
rect 1548 11651 1554 11654
rect 156 11614 162 11617
rect 126 11608 162 11614
rect 810 11614 816 11617
rect 810 11608 1584 11614
rect 126 11574 138 11608
rect 1572 11574 1584 11608
rect 126 11568 162 11574
rect 156 11565 162 11568
rect 810 11568 1584 11574
rect 810 11565 816 11568
rect 894 11528 900 11531
rect 126 11522 900 11528
rect 1548 11528 1554 11531
rect 1548 11522 1584 11528
rect 126 11488 138 11522
rect 1572 11488 1584 11522
rect 126 11482 900 11488
rect 894 11479 900 11482
rect 1548 11482 1584 11488
rect 1548 11479 1554 11482
rect 156 11442 162 11445
rect 126 11436 162 11442
rect 810 11442 816 11445
rect 810 11436 1584 11442
rect 126 11402 138 11436
rect 1572 11402 1584 11436
rect 126 11396 162 11402
rect 156 11393 162 11396
rect 810 11396 1584 11402
rect 810 11393 816 11396
rect 894 11356 900 11359
rect 126 11350 900 11356
rect 1548 11356 1554 11359
rect 1548 11350 1584 11356
rect 126 11316 138 11350
rect 1572 11316 1584 11350
rect 126 11310 900 11316
rect 894 11307 900 11310
rect 1548 11310 1584 11316
rect 1548 11307 1554 11310
rect 156 11270 162 11273
rect 126 11264 162 11270
rect 810 11270 816 11273
rect 810 11264 1584 11270
rect 126 11230 138 11264
rect 1572 11230 1584 11264
rect 126 11224 162 11230
rect 156 11221 162 11224
rect 810 11224 1584 11230
rect 810 11221 816 11224
rect 894 11184 900 11187
rect 126 11178 900 11184
rect 1548 11184 1554 11187
rect 1548 11178 1584 11184
rect 126 11144 138 11178
rect 1572 11144 1584 11178
rect 126 11138 900 11144
rect 894 11135 900 11138
rect 1548 11138 1584 11144
rect 1548 11135 1554 11138
rect 156 11098 162 11101
rect 126 11092 162 11098
rect 810 11098 816 11101
rect 810 11092 1584 11098
rect 126 11058 138 11092
rect 1572 11058 1584 11092
rect 126 11052 162 11058
rect 156 11049 162 11052
rect 810 11052 1584 11058
rect 810 11049 816 11052
rect 894 11012 900 11015
rect 126 11006 900 11012
rect 1548 11012 1554 11015
rect 1548 11006 1584 11012
rect 126 10972 138 11006
rect 1572 10972 1584 11006
rect 126 10966 900 10972
rect 894 10963 900 10966
rect 1548 10966 1584 10972
rect 1548 10963 1554 10966
rect 156 10926 162 10929
rect 126 10920 162 10926
rect 810 10926 816 10929
rect 810 10920 1584 10926
rect 126 10886 138 10920
rect 1572 10886 1584 10920
rect 126 10880 162 10886
rect 156 10877 162 10880
rect 810 10880 1584 10886
rect 810 10877 816 10880
rect 894 10840 900 10843
rect 126 10834 900 10840
rect 1548 10840 1554 10843
rect 1548 10834 1584 10840
rect 126 10800 138 10834
rect 1572 10800 1584 10834
rect 126 10794 900 10800
rect 894 10791 900 10794
rect 1548 10794 1584 10800
rect 1548 10791 1554 10794
rect 156 10754 162 10757
rect 126 10748 162 10754
rect 810 10754 816 10757
rect 810 10748 1584 10754
rect 126 10714 138 10748
rect 1572 10714 1584 10748
rect 126 10708 162 10714
rect 156 10705 162 10708
rect 810 10708 1584 10714
rect 810 10705 816 10708
rect 894 10668 900 10671
rect 126 10662 900 10668
rect 1548 10668 1554 10671
rect 1548 10662 1584 10668
rect 126 10628 138 10662
rect 1572 10628 1584 10662
rect 126 10622 900 10628
rect 894 10619 900 10622
rect 1548 10622 1584 10628
rect 1548 10619 1554 10622
rect 156 10582 162 10585
rect 126 10576 162 10582
rect 810 10582 816 10585
rect 810 10576 1584 10582
rect 126 10542 138 10576
rect 1572 10542 1584 10576
rect 126 10536 162 10542
rect 156 10533 162 10536
rect 810 10536 1584 10542
rect 810 10533 816 10536
rect 894 10496 900 10499
rect 126 10490 900 10496
rect 1548 10496 1554 10499
rect 1548 10490 1584 10496
rect 126 10456 138 10490
rect 1572 10456 1584 10490
rect 126 10450 900 10456
rect 894 10447 900 10450
rect 1548 10450 1584 10456
rect 1548 10447 1554 10450
rect 156 10410 162 10413
rect 126 10404 162 10410
rect 810 10410 816 10413
rect 810 10404 1584 10410
rect 126 10370 138 10404
rect 1572 10370 1584 10404
rect 126 10364 162 10370
rect 156 10361 162 10364
rect 810 10364 1584 10370
rect 810 10361 816 10364
rect 894 10324 900 10327
rect 126 10318 900 10324
rect 1548 10324 1554 10327
rect 1548 10318 1584 10324
rect 126 10284 138 10318
rect 1572 10284 1584 10318
rect 126 10278 900 10284
rect 894 10275 900 10278
rect 1548 10278 1584 10284
rect 1548 10275 1554 10278
rect 156 10238 162 10241
rect 126 10232 162 10238
rect 810 10238 816 10241
rect 810 10232 1584 10238
rect 126 10198 138 10232
rect 1572 10198 1584 10232
rect 126 10192 162 10198
rect 156 10189 162 10192
rect 810 10192 1584 10198
rect 810 10189 816 10192
rect 894 10152 900 10155
rect 126 10146 900 10152
rect 1548 10152 1554 10155
rect 1548 10146 1584 10152
rect 126 10112 138 10146
rect 1572 10112 1584 10146
rect 126 10106 900 10112
rect 894 10103 900 10106
rect 1548 10106 1584 10112
rect 1548 10103 1554 10106
rect 156 10066 162 10069
rect 126 10060 162 10066
rect 810 10066 816 10069
rect 810 10060 1584 10066
rect 126 10026 138 10060
rect 1572 10026 1584 10060
rect 126 10020 162 10026
rect 156 10017 162 10020
rect 810 10020 1584 10026
rect 810 10017 816 10020
rect 894 9980 900 9983
rect 126 9974 900 9980
rect 1548 9980 1554 9983
rect 1548 9974 1584 9980
rect 126 9940 138 9974
rect 1572 9940 1584 9974
rect 126 9934 900 9940
rect 894 9931 900 9934
rect 1548 9934 1584 9940
rect 1548 9931 1554 9934
rect 156 9894 162 9897
rect 126 9888 162 9894
rect 810 9894 816 9897
rect 810 9888 1584 9894
rect 126 9854 138 9888
rect 1572 9854 1584 9888
rect 126 9848 162 9854
rect 156 9845 162 9848
rect 810 9848 1584 9854
rect 810 9845 816 9848
rect 894 9808 900 9811
rect 126 9802 900 9808
rect 1548 9808 1554 9811
rect 1548 9802 1584 9808
rect 126 9768 138 9802
rect 1572 9768 1584 9802
rect 126 9762 900 9768
rect 894 9759 900 9762
rect 1548 9762 1584 9768
rect 1548 9759 1554 9762
rect 156 9722 162 9725
rect 126 9716 162 9722
rect 810 9722 816 9725
rect 810 9716 1584 9722
rect 126 9682 138 9716
rect 1572 9682 1584 9716
rect 126 9676 162 9682
rect 156 9673 162 9676
rect 810 9676 1584 9682
rect 810 9673 816 9676
rect 894 9636 900 9639
rect 126 9630 900 9636
rect 1548 9636 1554 9639
rect 1548 9630 1584 9636
rect 126 9596 138 9630
rect 1572 9596 1584 9630
rect 126 9590 900 9596
rect 894 9587 900 9590
rect 1548 9590 1584 9596
rect 1548 9587 1554 9590
rect 156 9550 162 9553
rect 126 9544 162 9550
rect 810 9550 816 9553
rect 810 9544 1584 9550
rect 126 9510 138 9544
rect 1572 9510 1584 9544
rect 126 9504 162 9510
rect 156 9501 162 9504
rect 810 9504 1584 9510
rect 810 9501 816 9504
rect 894 9464 900 9467
rect 126 9458 900 9464
rect 1548 9464 1554 9467
rect 1548 9458 1584 9464
rect 126 9424 138 9458
rect 1572 9424 1584 9458
rect 126 9418 900 9424
rect 894 9415 900 9418
rect 1548 9418 1584 9424
rect 1548 9415 1554 9418
rect 156 9378 162 9381
rect 126 9372 162 9378
rect 810 9378 816 9381
rect 810 9372 1584 9378
rect 126 9338 138 9372
rect 1572 9338 1584 9372
rect 126 9332 162 9338
rect 156 9329 162 9332
rect 810 9332 1584 9338
rect 810 9329 816 9332
rect 894 9292 900 9295
rect 126 9286 900 9292
rect 1548 9292 1554 9295
rect 1548 9286 1584 9292
rect 126 9252 138 9286
rect 1572 9252 1584 9286
rect 126 9246 900 9252
rect 894 9243 900 9246
rect 1548 9246 1584 9252
rect 1548 9243 1554 9246
rect 156 9206 162 9209
rect 126 9200 162 9206
rect 810 9206 816 9209
rect 810 9200 1584 9206
rect 126 9166 138 9200
rect 1572 9166 1584 9200
rect 126 9160 162 9166
rect 156 9157 162 9160
rect 810 9160 1584 9166
rect 810 9157 816 9160
rect 894 9120 900 9123
rect 126 9114 900 9120
rect 1548 9120 1554 9123
rect 1548 9114 1584 9120
rect 126 9080 138 9114
rect 1572 9080 1584 9114
rect 126 9074 900 9080
rect 894 9071 900 9074
rect 1548 9074 1584 9080
rect 1548 9071 1554 9074
rect 156 9034 162 9037
rect 126 9028 162 9034
rect 810 9034 816 9037
rect 810 9028 1584 9034
rect 126 8994 138 9028
rect 1572 8994 1584 9028
rect 126 8988 162 8994
rect 156 8985 162 8988
rect 810 8988 1584 8994
rect 810 8985 816 8988
rect 894 8948 900 8951
rect 126 8942 900 8948
rect 1548 8948 1554 8951
rect 1548 8942 1584 8948
rect 126 8908 138 8942
rect 1572 8908 1584 8942
rect 126 8902 900 8908
rect 894 8899 900 8902
rect 1548 8902 1584 8908
rect 1548 8899 1554 8902
rect 156 8862 162 8865
rect 126 8856 162 8862
rect 810 8862 816 8865
rect 810 8856 1584 8862
rect 126 8822 138 8856
rect 1572 8822 1584 8856
rect 126 8816 162 8822
rect 156 8813 162 8816
rect 810 8816 1584 8822
rect 810 8813 816 8816
rect 894 8776 900 8779
rect 126 8770 900 8776
rect 1548 8776 1554 8779
rect 1548 8770 1584 8776
rect 126 8736 138 8770
rect 1572 8736 1584 8770
rect 126 8730 900 8736
rect 894 8727 900 8730
rect 1548 8730 1584 8736
rect 1548 8727 1554 8730
rect 156 8690 162 8693
rect 126 8684 162 8690
rect 810 8690 816 8693
rect 810 8684 1584 8690
rect 126 8650 138 8684
rect 1572 8650 1584 8684
rect 126 8644 162 8650
rect 156 8641 162 8644
rect 810 8644 1584 8650
rect 810 8641 816 8644
rect 894 8604 900 8607
rect 126 8598 900 8604
rect 1548 8604 1554 8607
rect 1548 8598 1584 8604
rect 126 8564 138 8598
rect 1572 8564 1584 8598
rect 126 8558 900 8564
rect 894 8555 900 8558
rect 1548 8558 1584 8564
rect 1548 8555 1554 8558
rect 156 8518 162 8521
rect 126 8512 162 8518
rect 810 8518 816 8521
rect 810 8512 1584 8518
rect 126 8478 138 8512
rect 1572 8478 1584 8512
rect 126 8472 162 8478
rect 156 8469 162 8472
rect 810 8472 1584 8478
rect 810 8469 816 8472
rect 894 8432 900 8435
rect 126 8426 900 8432
rect 1548 8432 1554 8435
rect 1548 8426 1584 8432
rect 126 8392 138 8426
rect 1572 8392 1584 8426
rect 126 8386 900 8392
rect 894 8383 900 8386
rect 1548 8386 1584 8392
rect 1548 8383 1554 8386
rect 156 8346 162 8349
rect 126 8340 162 8346
rect 810 8346 816 8349
rect 810 8340 1584 8346
rect 126 8306 138 8340
rect 1572 8306 1584 8340
rect 126 8300 162 8306
rect 156 8297 162 8300
rect 810 8300 1584 8306
rect 810 8297 816 8300
rect 894 8260 900 8263
rect 126 8254 900 8260
rect 1548 8260 1554 8263
rect 1548 8254 1584 8260
rect 126 8220 138 8254
rect 1572 8220 1584 8254
rect 126 8214 900 8220
rect 894 8211 900 8214
rect 1548 8214 1584 8220
rect 1548 8211 1554 8214
rect 156 8174 162 8177
rect 126 8168 162 8174
rect 810 8174 816 8177
rect 810 8168 1584 8174
rect 126 8134 138 8168
rect 1572 8134 1584 8168
rect 126 8128 162 8134
rect 156 8125 162 8128
rect 810 8128 1584 8134
rect 810 8125 816 8128
rect 894 8088 900 8091
rect 126 8082 900 8088
rect 1548 8088 1554 8091
rect 1548 8082 1584 8088
rect 126 8048 138 8082
rect 1572 8048 1584 8082
rect 126 8042 900 8048
rect 894 8039 900 8042
rect 1548 8042 1584 8048
rect 1548 8039 1554 8042
rect 156 8002 162 8005
rect 126 7996 162 8002
rect 810 8002 816 8005
rect 810 7996 1584 8002
rect 126 7962 138 7996
rect 1572 7962 1584 7996
rect 126 7956 162 7962
rect 156 7953 162 7956
rect 810 7956 1584 7962
rect 810 7953 816 7956
rect 894 7916 900 7919
rect 126 7910 900 7916
rect 1548 7916 1554 7919
rect 1548 7910 1584 7916
rect 126 7876 138 7910
rect 1572 7876 1584 7910
rect 126 7870 900 7876
rect 894 7867 900 7870
rect 1548 7870 1584 7876
rect 1548 7867 1554 7870
rect 156 7830 162 7833
rect 126 7824 162 7830
rect 810 7830 816 7833
rect 810 7824 1584 7830
rect 126 7790 138 7824
rect 1572 7790 1584 7824
rect 126 7784 162 7790
rect 156 7781 162 7784
rect 810 7784 1584 7790
rect 810 7781 816 7784
rect 894 7744 900 7747
rect 126 7738 900 7744
rect 1548 7744 1554 7747
rect 1548 7738 1584 7744
rect 126 7704 138 7738
rect 1572 7704 1584 7738
rect 126 7698 900 7704
rect 894 7695 900 7698
rect 1548 7698 1584 7704
rect 1548 7695 1554 7698
rect 156 7658 162 7661
rect 126 7652 162 7658
rect 810 7658 816 7661
rect 810 7652 1584 7658
rect 126 7618 138 7652
rect 1572 7618 1584 7652
rect 126 7612 162 7618
rect 156 7609 162 7612
rect 810 7612 1584 7618
rect 810 7609 816 7612
rect 894 7572 900 7575
rect 126 7566 900 7572
rect 1548 7572 1554 7575
rect 1548 7566 1584 7572
rect 126 7532 138 7566
rect 1572 7532 1584 7566
rect 126 7526 900 7532
rect 894 7523 900 7526
rect 1548 7526 1584 7532
rect 1548 7523 1554 7526
rect 156 7486 162 7489
rect 126 7480 162 7486
rect 810 7486 816 7489
rect 810 7480 1584 7486
rect 126 7446 138 7480
rect 1572 7446 1584 7480
rect 126 7440 162 7446
rect 156 7437 162 7440
rect 810 7440 1584 7446
rect 810 7437 816 7440
rect 894 7400 900 7403
rect 126 7394 900 7400
rect 1548 7400 1554 7403
rect 1548 7394 1584 7400
rect 126 7360 138 7394
rect 1572 7360 1584 7394
rect 126 7354 900 7360
rect 894 7351 900 7354
rect 1548 7354 1584 7360
rect 1548 7351 1554 7354
rect 156 7314 162 7317
rect 126 7308 162 7314
rect 810 7314 816 7317
rect 810 7308 1584 7314
rect 126 7274 138 7308
rect 1572 7274 1584 7308
rect 126 7268 162 7274
rect 156 7265 162 7268
rect 810 7268 1584 7274
rect 810 7265 816 7268
rect 894 7228 900 7231
rect 126 7222 900 7228
rect 1548 7228 1554 7231
rect 1548 7222 1584 7228
rect 126 7188 138 7222
rect 1572 7188 1584 7222
rect 126 7182 900 7188
rect 894 7179 900 7182
rect 1548 7182 1584 7188
rect 1548 7179 1554 7182
rect 156 7142 162 7145
rect 126 7136 162 7142
rect 810 7142 816 7145
rect 810 7136 1584 7142
rect 126 7102 138 7136
rect 1572 7102 1584 7136
rect 126 7096 162 7102
rect 156 7093 162 7096
rect 810 7096 1584 7102
rect 810 7093 816 7096
rect 894 7056 900 7059
rect 126 7050 900 7056
rect 1548 7056 1554 7059
rect 1548 7050 1584 7056
rect 126 7016 138 7050
rect 1572 7016 1584 7050
rect 126 7010 900 7016
rect 894 7007 900 7010
rect 1548 7010 1584 7016
rect 1548 7007 1554 7010
rect 156 6970 162 6973
rect 126 6964 162 6970
rect 810 6970 816 6973
rect 810 6964 1584 6970
rect 126 6930 138 6964
rect 1572 6930 1584 6964
rect 126 6924 162 6930
rect 156 6921 162 6924
rect 810 6924 1584 6930
rect 810 6921 816 6924
rect 894 6884 900 6887
rect 126 6878 900 6884
rect 1548 6884 1554 6887
rect 1548 6878 1584 6884
rect 126 6844 138 6878
rect 1572 6844 1584 6878
rect 126 6838 900 6844
rect 894 6835 900 6838
rect 1548 6838 1584 6844
rect 1548 6835 1554 6838
rect 156 6798 162 6801
rect 126 6792 162 6798
rect 810 6798 816 6801
rect 810 6792 1584 6798
rect 126 6758 138 6792
rect 1572 6758 1584 6792
rect 126 6752 162 6758
rect 156 6749 162 6752
rect 810 6752 1584 6758
rect 810 6749 816 6752
rect 894 6712 900 6715
rect 126 6706 900 6712
rect 1548 6712 1554 6715
rect 1548 6706 1584 6712
rect 126 6672 138 6706
rect 1572 6672 1584 6706
rect 126 6666 900 6672
rect 894 6663 900 6666
rect 1548 6666 1584 6672
rect 1548 6663 1554 6666
rect 156 6626 162 6629
rect 126 6620 162 6626
rect 810 6626 816 6629
rect 810 6620 1584 6626
rect 126 6586 138 6620
rect 1572 6586 1584 6620
rect 126 6580 162 6586
rect 156 6577 162 6580
rect 810 6580 1584 6586
rect 810 6577 816 6580
rect 894 6540 900 6543
rect 126 6534 900 6540
rect 1548 6540 1554 6543
rect 1548 6534 1584 6540
rect 126 6500 138 6534
rect 1572 6500 1584 6534
rect 126 6494 900 6500
rect 894 6491 900 6494
rect 1548 6494 1584 6500
rect 1548 6491 1554 6494
rect 156 6454 162 6457
rect 126 6448 162 6454
rect 810 6454 816 6457
rect 810 6448 1584 6454
rect 126 6414 138 6448
rect 1572 6414 1584 6448
rect 126 6408 162 6414
rect 156 6405 162 6408
rect 810 6408 1584 6414
rect 810 6405 816 6408
rect 894 6368 900 6371
rect 126 6362 900 6368
rect 1548 6368 1554 6371
rect 1548 6362 1584 6368
rect 126 6328 138 6362
rect 1572 6328 1584 6362
rect 126 6322 900 6328
rect 894 6319 900 6322
rect 1548 6322 1584 6328
rect 1548 6319 1554 6322
rect 156 6282 162 6285
rect 126 6276 162 6282
rect 810 6282 816 6285
rect 810 6276 1584 6282
rect 126 6242 138 6276
rect 1572 6242 1584 6276
rect 126 6236 162 6242
rect 156 6233 162 6236
rect 810 6236 1584 6242
rect 810 6233 816 6236
rect 894 6196 900 6199
rect 126 6190 900 6196
rect 1548 6196 1554 6199
rect 1548 6190 1584 6196
rect 126 6156 138 6190
rect 1572 6156 1584 6190
rect 126 6150 900 6156
rect 894 6147 900 6150
rect 1548 6150 1584 6156
rect 1548 6147 1554 6150
rect 156 6110 162 6113
rect 126 6104 162 6110
rect 810 6110 816 6113
rect 810 6104 1584 6110
rect 126 6070 138 6104
rect 1572 6070 1584 6104
rect 126 6064 162 6070
rect 156 6061 162 6064
rect 810 6064 1584 6070
rect 810 6061 816 6064
rect 894 6024 900 6027
rect 126 6018 900 6024
rect 1548 6024 1554 6027
rect 1548 6018 1584 6024
rect 126 5984 138 6018
rect 1572 5984 1584 6018
rect 126 5978 900 5984
rect 894 5975 900 5978
rect 1548 5978 1584 5984
rect 1548 5975 1554 5978
rect 156 5938 162 5941
rect 126 5932 162 5938
rect 810 5938 816 5941
rect 810 5932 1584 5938
rect 126 5898 138 5932
rect 1572 5898 1584 5932
rect 126 5892 162 5898
rect 156 5889 162 5892
rect 810 5892 1584 5898
rect 810 5889 816 5892
rect 894 5852 900 5855
rect 126 5846 900 5852
rect 1548 5852 1554 5855
rect 1548 5846 1584 5852
rect 126 5812 138 5846
rect 1572 5812 1584 5846
rect 126 5806 900 5812
rect 894 5803 900 5806
rect 1548 5806 1584 5812
rect 1548 5803 1554 5806
rect 156 5766 162 5769
rect 126 5760 162 5766
rect 810 5766 816 5769
rect 810 5760 1584 5766
rect 126 5726 138 5760
rect 1572 5726 1584 5760
rect 126 5720 162 5726
rect 156 5717 162 5720
rect 810 5720 1584 5726
rect 810 5717 816 5720
rect 894 5680 900 5683
rect 126 5674 900 5680
rect 1548 5680 1554 5683
rect 1548 5674 1584 5680
rect 126 5640 138 5674
rect 1572 5640 1584 5674
rect 126 5634 900 5640
rect 894 5631 900 5634
rect 1548 5634 1584 5640
rect 1548 5631 1554 5634
rect 156 5594 162 5597
rect 126 5588 162 5594
rect 810 5594 816 5597
rect 810 5588 1584 5594
rect 126 5554 138 5588
rect 1572 5554 1584 5588
rect 126 5548 162 5554
rect 156 5545 162 5548
rect 810 5548 1584 5554
rect 810 5545 816 5548
rect 894 5508 900 5511
rect 126 5502 900 5508
rect 1548 5508 1554 5511
rect 1548 5502 1584 5508
rect 126 5468 138 5502
rect 1572 5468 1584 5502
rect 126 5462 900 5468
rect 894 5459 900 5462
rect 1548 5462 1584 5468
rect 1548 5459 1554 5462
rect 156 5422 162 5425
rect 126 5416 162 5422
rect 810 5422 816 5425
rect 810 5416 1584 5422
rect 126 5382 138 5416
rect 1572 5382 1584 5416
rect 126 5376 162 5382
rect 156 5373 162 5376
rect 810 5376 1584 5382
rect 810 5373 816 5376
rect 894 5336 900 5339
rect 126 5330 900 5336
rect 1548 5336 1554 5339
rect 1548 5330 1584 5336
rect 126 5296 138 5330
rect 1572 5296 1584 5330
rect 126 5290 900 5296
rect 894 5287 900 5290
rect 1548 5290 1584 5296
rect 1548 5287 1554 5290
rect 156 5250 162 5253
rect 126 5244 162 5250
rect 810 5250 816 5253
rect 810 5244 1584 5250
rect 126 5210 138 5244
rect 1572 5210 1584 5244
rect 126 5204 162 5210
rect 156 5201 162 5204
rect 810 5204 1584 5210
rect 810 5201 816 5204
rect 894 5164 900 5167
rect 126 5158 900 5164
rect 1548 5164 1554 5167
rect 1548 5158 1584 5164
rect 126 5124 138 5158
rect 1572 5124 1584 5158
rect 126 5118 900 5124
rect 894 5115 900 5118
rect 1548 5118 1584 5124
rect 1548 5115 1554 5118
rect 156 5078 162 5081
rect 126 5072 162 5078
rect 810 5078 816 5081
rect 810 5072 1584 5078
rect 126 5038 138 5072
rect 1572 5038 1584 5072
rect 126 5032 162 5038
rect 156 5029 162 5032
rect 810 5032 1584 5038
rect 810 5029 816 5032
rect 894 4992 900 4995
rect 126 4986 900 4992
rect 1548 4992 1554 4995
rect 1548 4986 1584 4992
rect 126 4952 138 4986
rect 1572 4952 1584 4986
rect 126 4946 900 4952
rect 894 4943 900 4946
rect 1548 4946 1584 4952
rect 1548 4943 1554 4946
rect 156 4906 162 4909
rect 126 4900 162 4906
rect 810 4906 816 4909
rect 810 4900 1584 4906
rect 126 4866 138 4900
rect 1572 4866 1584 4900
rect 126 4860 162 4866
rect 156 4857 162 4860
rect 810 4860 1584 4866
rect 810 4857 816 4860
rect 894 4820 900 4823
rect 126 4814 900 4820
rect 1548 4820 1554 4823
rect 1548 4814 1584 4820
rect 126 4780 138 4814
rect 1572 4780 1584 4814
rect 126 4774 900 4780
rect 894 4771 900 4774
rect 1548 4774 1584 4780
rect 1548 4771 1554 4774
rect 156 4734 162 4737
rect 126 4728 162 4734
rect 810 4734 816 4737
rect 810 4728 1584 4734
rect 126 4694 138 4728
rect 1572 4694 1584 4728
rect 126 4688 162 4694
rect 156 4685 162 4688
rect 810 4688 1584 4694
rect 810 4685 816 4688
rect 894 4648 900 4651
rect 126 4642 900 4648
rect 1548 4648 1554 4651
rect 1548 4642 1584 4648
rect 126 4608 138 4642
rect 1572 4608 1584 4642
rect 126 4602 900 4608
rect 894 4599 900 4602
rect 1548 4602 1584 4608
rect 1548 4599 1554 4602
rect 156 4562 162 4565
rect 126 4556 162 4562
rect 810 4562 816 4565
rect 810 4556 1584 4562
rect 126 4522 138 4556
rect 1572 4522 1584 4556
rect 126 4516 162 4522
rect 156 4513 162 4516
rect 810 4516 1584 4522
rect 810 4513 816 4516
rect 894 4476 900 4479
rect 126 4470 900 4476
rect 1548 4476 1554 4479
rect 1548 4470 1584 4476
rect 126 4436 138 4470
rect 1572 4436 1584 4470
rect 126 4430 900 4436
rect 894 4427 900 4430
rect 1548 4430 1584 4436
rect 1548 4427 1554 4430
rect 156 4390 162 4393
rect 126 4384 162 4390
rect 810 4390 816 4393
rect 810 4384 1584 4390
rect 126 4350 138 4384
rect 1572 4350 1584 4384
rect 126 4344 162 4350
rect 156 4341 162 4344
rect 810 4344 1584 4350
rect 810 4341 816 4344
rect 894 4304 900 4307
rect 126 4298 900 4304
rect 1548 4304 1554 4307
rect 1548 4298 1584 4304
rect 126 4264 138 4298
rect 1572 4264 1584 4298
rect 126 4258 900 4264
rect 894 4255 900 4258
rect 1548 4258 1584 4264
rect 1548 4255 1554 4258
rect 156 4218 162 4221
rect 126 4212 162 4218
rect 810 4218 816 4221
rect 810 4212 1584 4218
rect 126 4178 138 4212
rect 1572 4178 1584 4212
rect 126 4172 162 4178
rect 156 4169 162 4172
rect 810 4172 1584 4178
rect 810 4169 816 4172
rect 894 4132 900 4135
rect 126 4126 900 4132
rect 1548 4132 1554 4135
rect 1548 4126 1584 4132
rect 126 4092 138 4126
rect 1572 4092 1584 4126
rect 126 4086 900 4092
rect 894 4083 900 4086
rect 1548 4086 1584 4092
rect 1548 4083 1554 4086
rect 156 4046 162 4049
rect 126 4040 162 4046
rect 810 4046 816 4049
rect 810 4040 1584 4046
rect 126 4006 138 4040
rect 1572 4006 1584 4040
rect 126 4000 162 4006
rect 156 3997 162 4000
rect 810 4000 1584 4006
rect 810 3997 816 4000
rect 894 3960 900 3963
rect 126 3954 900 3960
rect 1548 3960 1554 3963
rect 1548 3954 1584 3960
rect 126 3920 138 3954
rect 1572 3920 1584 3954
rect 126 3914 900 3920
rect 894 3911 900 3914
rect 1548 3914 1584 3920
rect 1548 3911 1554 3914
rect 156 3874 162 3877
rect 126 3868 162 3874
rect 810 3874 816 3877
rect 810 3868 1584 3874
rect 126 3834 138 3868
rect 1572 3834 1584 3868
rect 126 3828 162 3834
rect 156 3825 162 3828
rect 810 3828 1584 3834
rect 810 3825 816 3828
rect 894 3788 900 3791
rect 126 3782 900 3788
rect 1548 3788 1554 3791
rect 1548 3782 1584 3788
rect 126 3748 138 3782
rect 1572 3748 1584 3782
rect 126 3742 900 3748
rect 894 3739 900 3742
rect 1548 3742 1584 3748
rect 1548 3739 1554 3742
rect 156 3702 162 3705
rect 126 3696 162 3702
rect 810 3702 816 3705
rect 810 3696 1584 3702
rect 126 3662 138 3696
rect 1572 3662 1584 3696
rect 126 3656 162 3662
rect 156 3653 162 3656
rect 810 3656 1584 3662
rect 810 3653 816 3656
rect 894 3616 900 3619
rect 126 3610 900 3616
rect 1548 3616 1554 3619
rect 1548 3610 1584 3616
rect 126 3576 138 3610
rect 1572 3576 1584 3610
rect 126 3570 900 3576
rect 894 3567 900 3570
rect 1548 3570 1584 3576
rect 1548 3567 1554 3570
rect 156 3530 162 3533
rect 126 3524 162 3530
rect 810 3530 816 3533
rect 810 3524 1584 3530
rect 126 3490 138 3524
rect 1572 3490 1584 3524
rect 126 3484 162 3490
rect 156 3481 162 3484
rect 810 3484 1584 3490
rect 810 3481 816 3484
rect 894 3444 900 3447
rect 126 3438 900 3444
rect 1548 3444 1554 3447
rect 1548 3438 1584 3444
rect 126 3404 138 3438
rect 1572 3404 1584 3438
rect 126 3398 900 3404
rect 894 3395 900 3398
rect 1548 3398 1584 3404
rect 1548 3395 1554 3398
rect 156 3358 162 3361
rect 126 3352 162 3358
rect 810 3358 816 3361
rect 810 3352 1584 3358
rect 126 3318 138 3352
rect 1572 3318 1584 3352
rect 126 3312 162 3318
rect 156 3309 162 3312
rect 810 3312 1584 3318
rect 810 3309 816 3312
rect 894 3272 900 3275
rect 126 3266 900 3272
rect 1548 3272 1554 3275
rect 1548 3266 1584 3272
rect 126 3232 138 3266
rect 1572 3232 1584 3266
rect 126 3226 900 3232
rect 894 3223 900 3226
rect 1548 3226 1584 3232
rect 1548 3223 1554 3226
rect 156 3186 162 3189
rect 126 3180 162 3186
rect 810 3186 816 3189
rect 810 3180 1584 3186
rect 126 3146 138 3180
rect 1572 3146 1584 3180
rect 126 3140 162 3146
rect 156 3137 162 3140
rect 810 3140 1584 3146
rect 810 3137 816 3140
rect 894 3100 900 3103
rect 126 3094 900 3100
rect 1548 3100 1554 3103
rect 1548 3094 1584 3100
rect 126 3060 138 3094
rect 1572 3060 1584 3094
rect 126 3054 900 3060
rect 894 3051 900 3054
rect 1548 3054 1584 3060
rect 1548 3051 1554 3054
rect 156 3014 162 3017
rect 126 3008 162 3014
rect 810 3014 816 3017
rect 810 3008 1584 3014
rect 126 2974 138 3008
rect 1572 2974 1584 3008
rect 126 2968 162 2974
rect 156 2965 162 2968
rect 810 2968 1584 2974
rect 810 2965 816 2968
rect 894 2928 900 2931
rect 126 2922 900 2928
rect 1548 2928 1554 2931
rect 1548 2922 1584 2928
rect 126 2888 138 2922
rect 1572 2888 1584 2922
rect 126 2882 900 2888
rect 894 2879 900 2882
rect 1548 2882 1584 2888
rect 1548 2879 1554 2882
rect 156 2842 162 2845
rect 126 2836 162 2842
rect 810 2842 816 2845
rect 810 2836 1584 2842
rect 126 2802 138 2836
rect 1572 2802 1584 2836
rect 126 2796 162 2802
rect 156 2793 162 2796
rect 810 2796 1584 2802
rect 810 2793 816 2796
rect 894 2756 900 2759
rect 126 2750 900 2756
rect 1548 2756 1554 2759
rect 1548 2750 1584 2756
rect 126 2716 138 2750
rect 1572 2716 1584 2750
rect 126 2710 900 2716
rect 894 2707 900 2710
rect 1548 2710 1584 2716
rect 1548 2707 1554 2710
rect 156 2670 162 2673
rect 126 2664 162 2670
rect 810 2670 816 2673
rect 810 2664 1584 2670
rect 126 2630 138 2664
rect 1572 2630 1584 2664
rect 126 2624 162 2630
rect 156 2621 162 2624
rect 810 2624 1584 2630
rect 810 2621 816 2624
rect 894 2584 900 2587
rect 126 2578 900 2584
rect 1548 2584 1554 2587
rect 1548 2578 1584 2584
rect 126 2544 138 2578
rect 1572 2544 1584 2578
rect 126 2538 900 2544
rect 894 2535 900 2538
rect 1548 2538 1584 2544
rect 1548 2535 1554 2538
rect 156 2498 162 2501
rect 126 2492 162 2498
rect 810 2498 816 2501
rect 810 2492 1584 2498
rect 126 2458 138 2492
rect 1572 2458 1584 2492
rect 126 2452 162 2458
rect 156 2449 162 2452
rect 810 2452 1584 2458
rect 810 2449 816 2452
rect 894 2412 900 2415
rect 126 2406 900 2412
rect 1548 2412 1554 2415
rect 1548 2406 1584 2412
rect 126 2372 138 2406
rect 1572 2372 1584 2406
rect 126 2366 900 2372
rect 894 2363 900 2366
rect 1548 2366 1584 2372
rect 1548 2363 1554 2366
rect 156 2326 162 2329
rect 126 2320 162 2326
rect 810 2326 816 2329
rect 810 2320 1584 2326
rect 126 2286 138 2320
rect 1572 2286 1584 2320
rect 126 2280 162 2286
rect 156 2277 162 2280
rect 810 2280 1584 2286
rect 810 2277 816 2280
rect 894 2240 900 2243
rect 126 2234 900 2240
rect 1548 2240 1554 2243
rect 1548 2234 1584 2240
rect 126 2200 138 2234
rect 1572 2200 1584 2234
rect 126 2194 900 2200
rect 894 2191 900 2194
rect 1548 2194 1584 2200
rect 1548 2191 1554 2194
rect 156 2154 162 2157
rect 126 2148 162 2154
rect 810 2154 816 2157
rect 810 2148 1584 2154
rect 126 2114 138 2148
rect 1572 2114 1584 2148
rect 126 2108 162 2114
rect 156 2105 162 2108
rect 810 2108 1584 2114
rect 810 2105 816 2108
rect 894 2068 900 2071
rect 126 2062 900 2068
rect 1548 2068 1554 2071
rect 1548 2062 1584 2068
rect 126 2028 138 2062
rect 1572 2028 1584 2062
rect 126 2022 900 2028
rect 894 2019 900 2022
rect 1548 2022 1584 2028
rect 1548 2019 1554 2022
rect 156 1982 162 1985
rect 126 1976 162 1982
rect 810 1982 816 1985
rect 810 1976 1584 1982
rect 126 1942 138 1976
rect 1572 1942 1584 1976
rect 126 1936 162 1942
rect 156 1933 162 1936
rect 810 1936 1584 1942
rect 810 1933 816 1936
rect 894 1896 900 1899
rect 126 1890 900 1896
rect 1548 1896 1554 1899
rect 1548 1890 1584 1896
rect 126 1856 138 1890
rect 1572 1856 1584 1890
rect 126 1850 900 1856
rect 894 1847 900 1850
rect 1548 1850 1584 1856
rect 1548 1847 1554 1850
rect 156 1810 162 1813
rect 126 1804 162 1810
rect 810 1810 816 1813
rect 810 1804 1584 1810
rect 126 1770 138 1804
rect 1572 1770 1584 1804
rect 126 1764 162 1770
rect 156 1761 162 1764
rect 810 1764 1584 1770
rect 810 1761 816 1764
rect 894 1724 900 1727
rect 126 1718 900 1724
rect 1548 1724 1554 1727
rect 1548 1718 1584 1724
rect 126 1684 138 1718
rect 1572 1684 1584 1718
rect 126 1678 900 1684
rect 894 1675 900 1678
rect 1548 1678 1584 1684
rect 1548 1675 1554 1678
rect 156 1638 162 1641
rect 126 1632 162 1638
rect 810 1638 816 1641
rect 810 1632 1584 1638
rect 126 1598 138 1632
rect 1572 1598 1584 1632
rect 126 1592 162 1598
rect 156 1589 162 1592
rect 810 1592 1584 1598
rect 810 1589 816 1592
rect 894 1552 900 1555
rect 126 1546 900 1552
rect 1548 1552 1554 1555
rect 1548 1546 1584 1552
rect 126 1512 138 1546
rect 1572 1512 1584 1546
rect 126 1506 900 1512
rect 894 1503 900 1506
rect 1548 1506 1584 1512
rect 1548 1503 1554 1506
rect 156 1466 162 1469
rect 126 1460 162 1466
rect 810 1466 816 1469
rect 810 1460 1584 1466
rect 126 1426 138 1460
rect 1572 1426 1584 1460
rect 126 1420 162 1426
rect 156 1417 162 1420
rect 810 1420 1584 1426
rect 810 1417 816 1420
rect 894 1380 900 1383
rect 126 1374 900 1380
rect 1548 1380 1554 1383
rect 1548 1374 1584 1380
rect 126 1340 138 1374
rect 1572 1340 1584 1374
rect 126 1334 900 1340
rect 894 1331 900 1334
rect 1548 1334 1584 1340
rect 1548 1331 1554 1334
rect 156 1294 162 1297
rect 126 1288 162 1294
rect 810 1294 816 1297
rect 810 1288 1584 1294
rect 126 1254 138 1288
rect 1572 1254 1584 1288
rect 126 1248 162 1254
rect 156 1245 162 1248
rect 810 1248 1584 1254
rect 810 1245 816 1248
rect 894 1208 900 1211
rect 126 1202 900 1208
rect 1548 1208 1554 1211
rect 1548 1202 1584 1208
rect 126 1168 138 1202
rect 1572 1168 1584 1202
rect 126 1162 900 1168
rect 894 1159 900 1162
rect 1548 1162 1584 1168
rect 1548 1159 1554 1162
rect 156 1122 162 1125
rect 126 1116 162 1122
rect 810 1122 816 1125
rect 810 1116 1584 1122
rect 126 1082 138 1116
rect 1572 1082 1584 1116
rect 126 1076 162 1082
rect 156 1073 162 1076
rect 810 1076 1584 1082
rect 810 1073 816 1076
rect 894 1036 900 1039
rect 126 1030 900 1036
rect 1548 1036 1554 1039
rect 1548 1030 1584 1036
rect 126 996 138 1030
rect 1572 996 1584 1030
rect 126 990 900 996
rect 894 987 900 990
rect 1548 990 1584 996
rect 1548 987 1554 990
rect 156 950 162 953
rect 126 944 162 950
rect 810 950 816 953
rect 810 944 1584 950
rect 126 910 138 944
rect 1572 910 1584 944
rect 126 904 162 910
rect 156 901 162 904
rect 810 904 1584 910
rect 810 901 816 904
rect 894 864 900 867
rect 126 858 900 864
rect 1548 864 1554 867
rect 1548 858 1584 864
rect 126 824 138 858
rect 1572 824 1584 858
rect 126 818 900 824
rect 894 815 900 818
rect 1548 818 1584 824
rect 1548 815 1554 818
rect 156 778 162 781
rect 126 772 162 778
rect 810 778 816 781
rect 810 772 1584 778
rect 126 738 138 772
rect 1572 738 1584 772
rect 126 732 162 738
rect 156 729 162 732
rect 810 732 1584 738
rect 810 729 816 732
rect 894 692 900 695
rect 126 686 900 692
rect 1548 692 1554 695
rect 1548 686 1584 692
rect 126 652 138 686
rect 1572 652 1584 686
rect 126 646 900 652
rect 894 643 900 646
rect 1548 646 1584 652
rect 1548 643 1554 646
rect 156 606 162 609
rect 126 600 162 606
rect 810 606 816 609
rect 810 600 1584 606
rect 126 566 138 600
rect 1572 566 1584 600
rect 126 560 162 566
rect 156 557 162 560
rect 810 560 1584 566
rect 810 557 816 560
rect 894 520 900 523
rect 126 514 900 520
rect 1548 520 1554 523
rect 1548 514 1584 520
rect 126 480 138 514
rect 1572 480 1584 514
rect 126 474 900 480
rect 894 471 900 474
rect 1548 474 1584 480
rect 1548 471 1554 474
rect 156 434 162 437
rect 126 428 162 434
rect 810 434 816 437
rect 810 428 1584 434
rect 126 394 138 428
rect 1572 394 1584 428
rect 126 388 162 394
rect 156 385 162 388
rect 810 388 1584 394
rect 810 385 816 388
rect 894 348 900 351
rect 126 342 900 348
rect 1548 348 1554 351
rect 1548 342 1584 348
rect 126 308 138 342
rect 1572 308 1584 342
rect 126 302 900 308
rect 894 299 900 302
rect 1548 302 1584 308
rect 1548 299 1554 302
rect 156 262 162 265
rect 126 256 162 262
rect 810 262 816 265
rect 810 256 1584 262
rect 126 222 138 256
rect 1572 222 1584 256
rect 126 216 162 222
rect 156 213 162 216
rect 810 216 1584 222
rect 810 213 816 216
rect 894 176 900 179
rect 126 170 900 176
rect 1548 176 1554 179
rect 1548 170 1584 176
rect 126 136 138 170
rect 1572 136 1584 170
rect 1618 163 1672 169
rect 126 130 900 136
rect 894 127 900 130
rect 1548 130 1584 136
rect 1548 127 1554 130
rect 30 76 76 100
rect 1704 100 1710 21190
rect 1744 100 1750 21190
rect 1704 76 1750 100
rect 30 70 1750 76
rect 30 36 100 70
rect 1680 36 1750 70
rect 30 30 1750 36
<< via1 >>
rect 900 21154 1548 21163
rect 900 21120 1548 21154
rect 900 21111 1548 21120
rect 1618 21111 1672 21121
rect 162 21068 810 21077
rect 162 21034 810 21068
rect 162 21025 810 21034
rect 900 20982 1548 20991
rect 900 20948 1548 20982
rect 900 20939 1548 20948
rect 162 20896 810 20905
rect 162 20862 810 20896
rect 162 20853 810 20862
rect 900 20810 1548 20819
rect 900 20776 1548 20810
rect 900 20767 1548 20776
rect 162 20724 810 20733
rect 162 20690 810 20724
rect 162 20681 810 20690
rect 900 20638 1548 20647
rect 900 20604 1548 20638
rect 900 20595 1548 20604
rect 162 20552 810 20561
rect 162 20518 810 20552
rect 162 20509 810 20518
rect 900 20466 1548 20475
rect 900 20432 1548 20466
rect 900 20423 1548 20432
rect 162 20380 810 20389
rect 162 20346 810 20380
rect 162 20337 810 20346
rect 900 20294 1548 20303
rect 900 20260 1548 20294
rect 900 20251 1548 20260
rect 162 20208 810 20217
rect 162 20174 810 20208
rect 162 20165 810 20174
rect 900 20122 1548 20131
rect 900 20088 1548 20122
rect 900 20079 1548 20088
rect 162 20036 810 20045
rect 162 20002 810 20036
rect 162 19993 810 20002
rect 900 19950 1548 19959
rect 900 19916 1548 19950
rect 900 19907 1548 19916
rect 162 19864 810 19873
rect 162 19830 810 19864
rect 162 19821 810 19830
rect 900 19778 1548 19787
rect 900 19744 1548 19778
rect 900 19735 1548 19744
rect 162 19692 810 19701
rect 162 19658 810 19692
rect 162 19649 810 19658
rect 900 19606 1548 19615
rect 900 19572 1548 19606
rect 900 19563 1548 19572
rect 162 19520 810 19529
rect 162 19486 810 19520
rect 162 19477 810 19486
rect 900 19434 1548 19443
rect 900 19400 1548 19434
rect 900 19391 1548 19400
rect 162 19348 810 19357
rect 162 19314 810 19348
rect 162 19305 810 19314
rect 900 19262 1548 19271
rect 900 19228 1548 19262
rect 900 19219 1548 19228
rect 162 19176 810 19185
rect 162 19142 810 19176
rect 162 19133 810 19142
rect 900 19090 1548 19099
rect 900 19056 1548 19090
rect 900 19047 1548 19056
rect 162 19004 810 19013
rect 162 18970 810 19004
rect 162 18961 810 18970
rect 900 18918 1548 18927
rect 900 18884 1548 18918
rect 900 18875 1548 18884
rect 162 18832 810 18841
rect 162 18798 810 18832
rect 162 18789 810 18798
rect 900 18746 1548 18755
rect 900 18712 1548 18746
rect 900 18703 1548 18712
rect 162 18660 810 18669
rect 162 18626 810 18660
rect 162 18617 810 18626
rect 900 18574 1548 18583
rect 900 18540 1548 18574
rect 900 18531 1548 18540
rect 162 18488 810 18497
rect 162 18454 810 18488
rect 162 18445 810 18454
rect 900 18402 1548 18411
rect 900 18368 1548 18402
rect 900 18359 1548 18368
rect 162 18316 810 18325
rect 162 18282 810 18316
rect 162 18273 810 18282
rect 900 18230 1548 18239
rect 900 18196 1548 18230
rect 900 18187 1548 18196
rect 162 18144 810 18153
rect 162 18110 810 18144
rect 162 18101 810 18110
rect 900 18058 1548 18067
rect 900 18024 1548 18058
rect 900 18015 1548 18024
rect 162 17972 810 17981
rect 162 17938 810 17972
rect 162 17929 810 17938
rect 900 17886 1548 17895
rect 900 17852 1548 17886
rect 900 17843 1548 17852
rect 162 17800 810 17809
rect 162 17766 810 17800
rect 162 17757 810 17766
rect 900 17714 1548 17723
rect 900 17680 1548 17714
rect 900 17671 1548 17680
rect 162 17628 810 17637
rect 162 17594 810 17628
rect 162 17585 810 17594
rect 900 17542 1548 17551
rect 900 17508 1548 17542
rect 900 17499 1548 17508
rect 162 17456 810 17465
rect 162 17422 810 17456
rect 162 17413 810 17422
rect 900 17370 1548 17379
rect 900 17336 1548 17370
rect 900 17327 1548 17336
rect 162 17284 810 17293
rect 162 17250 810 17284
rect 162 17241 810 17250
rect 900 17198 1548 17207
rect 900 17164 1548 17198
rect 900 17155 1548 17164
rect 162 17112 810 17121
rect 162 17078 810 17112
rect 162 17069 810 17078
rect 900 17026 1548 17035
rect 900 16992 1548 17026
rect 900 16983 1548 16992
rect 162 16940 810 16949
rect 162 16906 810 16940
rect 162 16897 810 16906
rect 900 16854 1548 16863
rect 900 16820 1548 16854
rect 900 16811 1548 16820
rect 162 16768 810 16777
rect 162 16734 810 16768
rect 162 16725 810 16734
rect 900 16682 1548 16691
rect 900 16648 1548 16682
rect 900 16639 1548 16648
rect 162 16596 810 16605
rect 162 16562 810 16596
rect 162 16553 810 16562
rect 900 16510 1548 16519
rect 900 16476 1548 16510
rect 900 16467 1548 16476
rect 162 16424 810 16433
rect 162 16390 810 16424
rect 162 16381 810 16390
rect 900 16338 1548 16347
rect 900 16304 1548 16338
rect 900 16295 1548 16304
rect 162 16252 810 16261
rect 162 16218 810 16252
rect 162 16209 810 16218
rect 900 16166 1548 16175
rect 900 16132 1548 16166
rect 900 16123 1548 16132
rect 162 16080 810 16089
rect 162 16046 810 16080
rect 162 16037 810 16046
rect 900 15994 1548 16003
rect 900 15960 1548 15994
rect 900 15951 1548 15960
rect 162 15908 810 15917
rect 162 15874 810 15908
rect 162 15865 810 15874
rect 900 15822 1548 15831
rect 900 15788 1548 15822
rect 900 15779 1548 15788
rect 162 15736 810 15745
rect 162 15702 810 15736
rect 162 15693 810 15702
rect 900 15650 1548 15659
rect 900 15616 1548 15650
rect 900 15607 1548 15616
rect 162 15564 810 15573
rect 162 15530 810 15564
rect 162 15521 810 15530
rect 900 15478 1548 15487
rect 900 15444 1548 15478
rect 900 15435 1548 15444
rect 162 15392 810 15401
rect 162 15358 810 15392
rect 162 15349 810 15358
rect 900 15306 1548 15315
rect 900 15272 1548 15306
rect 900 15263 1548 15272
rect 162 15220 810 15229
rect 162 15186 810 15220
rect 162 15177 810 15186
rect 900 15134 1548 15143
rect 900 15100 1548 15134
rect 900 15091 1548 15100
rect 162 15048 810 15057
rect 162 15014 810 15048
rect 162 15005 810 15014
rect 900 14962 1548 14971
rect 900 14928 1548 14962
rect 900 14919 1548 14928
rect 162 14876 810 14885
rect 162 14842 810 14876
rect 162 14833 810 14842
rect 900 14790 1548 14799
rect 900 14756 1548 14790
rect 900 14747 1548 14756
rect 162 14704 810 14713
rect 162 14670 810 14704
rect 162 14661 810 14670
rect 900 14618 1548 14627
rect 900 14584 1548 14618
rect 900 14575 1548 14584
rect 162 14532 810 14541
rect 162 14498 810 14532
rect 162 14489 810 14498
rect 900 14446 1548 14455
rect 900 14412 1548 14446
rect 900 14403 1548 14412
rect 162 14360 810 14369
rect 162 14326 810 14360
rect 162 14317 810 14326
rect 900 14274 1548 14283
rect 900 14240 1548 14274
rect 900 14231 1548 14240
rect 162 14188 810 14197
rect 162 14154 810 14188
rect 162 14145 810 14154
rect 900 14102 1548 14111
rect 900 14068 1548 14102
rect 900 14059 1548 14068
rect 162 14016 810 14025
rect 162 13982 810 14016
rect 162 13973 810 13982
rect 900 13930 1548 13939
rect 900 13896 1548 13930
rect 900 13887 1548 13896
rect 162 13844 810 13853
rect 162 13810 810 13844
rect 162 13801 810 13810
rect 900 13758 1548 13767
rect 900 13724 1548 13758
rect 900 13715 1548 13724
rect 162 13672 810 13681
rect 162 13638 810 13672
rect 162 13629 810 13638
rect 900 13586 1548 13595
rect 900 13552 1548 13586
rect 900 13543 1548 13552
rect 162 13500 810 13509
rect 162 13466 810 13500
rect 162 13457 810 13466
rect 900 13414 1548 13423
rect 900 13380 1548 13414
rect 900 13371 1548 13380
rect 162 13328 810 13337
rect 162 13294 810 13328
rect 162 13285 810 13294
rect 900 13242 1548 13251
rect 900 13208 1548 13242
rect 900 13199 1548 13208
rect 162 13156 810 13165
rect 162 13122 810 13156
rect 162 13113 810 13122
rect 900 13070 1548 13079
rect 900 13036 1548 13070
rect 900 13027 1548 13036
rect 162 12984 810 12993
rect 162 12950 810 12984
rect 162 12941 810 12950
rect 900 12898 1548 12907
rect 900 12864 1548 12898
rect 900 12855 1548 12864
rect 162 12812 810 12821
rect 162 12778 810 12812
rect 162 12769 810 12778
rect 900 12726 1548 12735
rect 900 12692 1548 12726
rect 900 12683 1548 12692
rect 162 12640 810 12649
rect 162 12606 810 12640
rect 162 12597 810 12606
rect 900 12554 1548 12563
rect 900 12520 1548 12554
rect 900 12511 1548 12520
rect 162 12468 810 12477
rect 162 12434 810 12468
rect 162 12425 810 12434
rect 900 12382 1548 12391
rect 900 12348 1548 12382
rect 900 12339 1548 12348
rect 162 12296 810 12305
rect 162 12262 810 12296
rect 162 12253 810 12262
rect 900 12210 1548 12219
rect 900 12176 1548 12210
rect 900 12167 1548 12176
rect 162 12124 810 12133
rect 162 12090 810 12124
rect 162 12081 810 12090
rect 900 12038 1548 12047
rect 900 12004 1548 12038
rect 900 11995 1548 12004
rect 162 11952 810 11961
rect 162 11918 810 11952
rect 162 11909 810 11918
rect 900 11866 1548 11875
rect 900 11832 1548 11866
rect 900 11823 1548 11832
rect 162 11780 810 11789
rect 162 11746 810 11780
rect 162 11737 810 11746
rect 900 11694 1548 11703
rect 900 11660 1548 11694
rect 900 11651 1548 11660
rect 162 11608 810 11617
rect 162 11574 810 11608
rect 162 11565 810 11574
rect 900 11522 1548 11531
rect 900 11488 1548 11522
rect 900 11479 1548 11488
rect 162 11436 810 11445
rect 162 11402 810 11436
rect 162 11393 810 11402
rect 900 11350 1548 11359
rect 900 11316 1548 11350
rect 900 11307 1548 11316
rect 162 11264 810 11273
rect 162 11230 810 11264
rect 162 11221 810 11230
rect 900 11178 1548 11187
rect 900 11144 1548 11178
rect 900 11135 1548 11144
rect 162 11092 810 11101
rect 162 11058 810 11092
rect 162 11049 810 11058
rect 900 11006 1548 11015
rect 900 10972 1548 11006
rect 900 10963 1548 10972
rect 162 10920 810 10929
rect 162 10886 810 10920
rect 162 10877 810 10886
rect 900 10834 1548 10843
rect 900 10800 1548 10834
rect 900 10791 1548 10800
rect 162 10748 810 10757
rect 162 10714 810 10748
rect 162 10705 810 10714
rect 900 10662 1548 10671
rect 900 10628 1548 10662
rect 900 10619 1548 10628
rect 162 10576 810 10585
rect 162 10542 810 10576
rect 162 10533 810 10542
rect 900 10490 1548 10499
rect 900 10456 1548 10490
rect 900 10447 1548 10456
rect 162 10404 810 10413
rect 162 10370 810 10404
rect 162 10361 810 10370
rect 900 10318 1548 10327
rect 900 10284 1548 10318
rect 900 10275 1548 10284
rect 162 10232 810 10241
rect 162 10198 810 10232
rect 162 10189 810 10198
rect 900 10146 1548 10155
rect 900 10112 1548 10146
rect 900 10103 1548 10112
rect 162 10060 810 10069
rect 162 10026 810 10060
rect 162 10017 810 10026
rect 900 9974 1548 9983
rect 900 9940 1548 9974
rect 900 9931 1548 9940
rect 162 9888 810 9897
rect 162 9854 810 9888
rect 162 9845 810 9854
rect 900 9802 1548 9811
rect 900 9768 1548 9802
rect 900 9759 1548 9768
rect 162 9716 810 9725
rect 162 9682 810 9716
rect 162 9673 810 9682
rect 900 9630 1548 9639
rect 900 9596 1548 9630
rect 900 9587 1548 9596
rect 162 9544 810 9553
rect 162 9510 810 9544
rect 162 9501 810 9510
rect 900 9458 1548 9467
rect 900 9424 1548 9458
rect 900 9415 1548 9424
rect 162 9372 810 9381
rect 162 9338 810 9372
rect 162 9329 810 9338
rect 900 9286 1548 9295
rect 900 9252 1548 9286
rect 900 9243 1548 9252
rect 162 9200 810 9209
rect 162 9166 810 9200
rect 162 9157 810 9166
rect 900 9114 1548 9123
rect 900 9080 1548 9114
rect 900 9071 1548 9080
rect 162 9028 810 9037
rect 162 8994 810 9028
rect 162 8985 810 8994
rect 900 8942 1548 8951
rect 900 8908 1548 8942
rect 900 8899 1548 8908
rect 162 8856 810 8865
rect 162 8822 810 8856
rect 162 8813 810 8822
rect 900 8770 1548 8779
rect 900 8736 1548 8770
rect 900 8727 1548 8736
rect 162 8684 810 8693
rect 162 8650 810 8684
rect 162 8641 810 8650
rect 900 8598 1548 8607
rect 900 8564 1548 8598
rect 900 8555 1548 8564
rect 162 8512 810 8521
rect 162 8478 810 8512
rect 162 8469 810 8478
rect 900 8426 1548 8435
rect 900 8392 1548 8426
rect 900 8383 1548 8392
rect 162 8340 810 8349
rect 162 8306 810 8340
rect 162 8297 810 8306
rect 900 8254 1548 8263
rect 900 8220 1548 8254
rect 900 8211 1548 8220
rect 162 8168 810 8177
rect 162 8134 810 8168
rect 162 8125 810 8134
rect 900 8082 1548 8091
rect 900 8048 1548 8082
rect 900 8039 1548 8048
rect 162 7996 810 8005
rect 162 7962 810 7996
rect 162 7953 810 7962
rect 900 7910 1548 7919
rect 900 7876 1548 7910
rect 900 7867 1548 7876
rect 162 7824 810 7833
rect 162 7790 810 7824
rect 162 7781 810 7790
rect 900 7738 1548 7747
rect 900 7704 1548 7738
rect 900 7695 1548 7704
rect 162 7652 810 7661
rect 162 7618 810 7652
rect 162 7609 810 7618
rect 900 7566 1548 7575
rect 900 7532 1548 7566
rect 900 7523 1548 7532
rect 162 7480 810 7489
rect 162 7446 810 7480
rect 162 7437 810 7446
rect 900 7394 1548 7403
rect 900 7360 1548 7394
rect 900 7351 1548 7360
rect 162 7308 810 7317
rect 162 7274 810 7308
rect 162 7265 810 7274
rect 900 7222 1548 7231
rect 900 7188 1548 7222
rect 900 7179 1548 7188
rect 162 7136 810 7145
rect 162 7102 810 7136
rect 162 7093 810 7102
rect 900 7050 1548 7059
rect 900 7016 1548 7050
rect 900 7007 1548 7016
rect 162 6964 810 6973
rect 162 6930 810 6964
rect 162 6921 810 6930
rect 900 6878 1548 6887
rect 900 6844 1548 6878
rect 900 6835 1548 6844
rect 162 6792 810 6801
rect 162 6758 810 6792
rect 162 6749 810 6758
rect 900 6706 1548 6715
rect 900 6672 1548 6706
rect 900 6663 1548 6672
rect 162 6620 810 6629
rect 162 6586 810 6620
rect 162 6577 810 6586
rect 900 6534 1548 6543
rect 900 6500 1548 6534
rect 900 6491 1548 6500
rect 162 6448 810 6457
rect 162 6414 810 6448
rect 162 6405 810 6414
rect 900 6362 1548 6371
rect 900 6328 1548 6362
rect 900 6319 1548 6328
rect 162 6276 810 6285
rect 162 6242 810 6276
rect 162 6233 810 6242
rect 900 6190 1548 6199
rect 900 6156 1548 6190
rect 900 6147 1548 6156
rect 162 6104 810 6113
rect 162 6070 810 6104
rect 162 6061 810 6070
rect 900 6018 1548 6027
rect 900 5984 1548 6018
rect 900 5975 1548 5984
rect 162 5932 810 5941
rect 162 5898 810 5932
rect 162 5889 810 5898
rect 900 5846 1548 5855
rect 900 5812 1548 5846
rect 900 5803 1548 5812
rect 162 5760 810 5769
rect 162 5726 810 5760
rect 162 5717 810 5726
rect 900 5674 1548 5683
rect 900 5640 1548 5674
rect 900 5631 1548 5640
rect 162 5588 810 5597
rect 162 5554 810 5588
rect 162 5545 810 5554
rect 900 5502 1548 5511
rect 900 5468 1548 5502
rect 900 5459 1548 5468
rect 162 5416 810 5425
rect 162 5382 810 5416
rect 162 5373 810 5382
rect 900 5330 1548 5339
rect 900 5296 1548 5330
rect 900 5287 1548 5296
rect 162 5244 810 5253
rect 162 5210 810 5244
rect 162 5201 810 5210
rect 900 5158 1548 5167
rect 900 5124 1548 5158
rect 900 5115 1548 5124
rect 162 5072 810 5081
rect 162 5038 810 5072
rect 162 5029 810 5038
rect 900 4986 1548 4995
rect 900 4952 1548 4986
rect 900 4943 1548 4952
rect 162 4900 810 4909
rect 162 4866 810 4900
rect 162 4857 810 4866
rect 900 4814 1548 4823
rect 900 4780 1548 4814
rect 900 4771 1548 4780
rect 162 4728 810 4737
rect 162 4694 810 4728
rect 162 4685 810 4694
rect 900 4642 1548 4651
rect 900 4608 1548 4642
rect 900 4599 1548 4608
rect 162 4556 810 4565
rect 162 4522 810 4556
rect 162 4513 810 4522
rect 900 4470 1548 4479
rect 900 4436 1548 4470
rect 900 4427 1548 4436
rect 162 4384 810 4393
rect 162 4350 810 4384
rect 162 4341 810 4350
rect 900 4298 1548 4307
rect 900 4264 1548 4298
rect 900 4255 1548 4264
rect 162 4212 810 4221
rect 162 4178 810 4212
rect 162 4169 810 4178
rect 900 4126 1548 4135
rect 900 4092 1548 4126
rect 900 4083 1548 4092
rect 162 4040 810 4049
rect 162 4006 810 4040
rect 162 3997 810 4006
rect 900 3954 1548 3963
rect 900 3920 1548 3954
rect 900 3911 1548 3920
rect 162 3868 810 3877
rect 162 3834 810 3868
rect 162 3825 810 3834
rect 900 3782 1548 3791
rect 900 3748 1548 3782
rect 900 3739 1548 3748
rect 162 3696 810 3705
rect 162 3662 810 3696
rect 162 3653 810 3662
rect 900 3610 1548 3619
rect 900 3576 1548 3610
rect 900 3567 1548 3576
rect 162 3524 810 3533
rect 162 3490 810 3524
rect 162 3481 810 3490
rect 900 3438 1548 3447
rect 900 3404 1548 3438
rect 900 3395 1548 3404
rect 162 3352 810 3361
rect 162 3318 810 3352
rect 162 3309 810 3318
rect 900 3266 1548 3275
rect 900 3232 1548 3266
rect 900 3223 1548 3232
rect 162 3180 810 3189
rect 162 3146 810 3180
rect 162 3137 810 3146
rect 900 3094 1548 3103
rect 900 3060 1548 3094
rect 900 3051 1548 3060
rect 162 3008 810 3017
rect 162 2974 810 3008
rect 162 2965 810 2974
rect 900 2922 1548 2931
rect 900 2888 1548 2922
rect 900 2879 1548 2888
rect 162 2836 810 2845
rect 162 2802 810 2836
rect 162 2793 810 2802
rect 900 2750 1548 2759
rect 900 2716 1548 2750
rect 900 2707 1548 2716
rect 162 2664 810 2673
rect 162 2630 810 2664
rect 162 2621 810 2630
rect 900 2578 1548 2587
rect 900 2544 1548 2578
rect 900 2535 1548 2544
rect 162 2492 810 2501
rect 162 2458 810 2492
rect 162 2449 810 2458
rect 900 2406 1548 2415
rect 900 2372 1548 2406
rect 900 2363 1548 2372
rect 162 2320 810 2329
rect 162 2286 810 2320
rect 162 2277 810 2286
rect 900 2234 1548 2243
rect 900 2200 1548 2234
rect 900 2191 1548 2200
rect 162 2148 810 2157
rect 162 2114 810 2148
rect 162 2105 810 2114
rect 900 2062 1548 2071
rect 900 2028 1548 2062
rect 900 2019 1548 2028
rect 162 1976 810 1985
rect 162 1942 810 1976
rect 162 1933 810 1942
rect 900 1890 1548 1899
rect 900 1856 1548 1890
rect 900 1847 1548 1856
rect 162 1804 810 1813
rect 162 1770 810 1804
rect 162 1761 810 1770
rect 900 1718 1548 1727
rect 900 1684 1548 1718
rect 900 1675 1548 1684
rect 162 1632 810 1641
rect 162 1598 810 1632
rect 162 1589 810 1598
rect 900 1546 1548 1555
rect 900 1512 1548 1546
rect 900 1503 1548 1512
rect 162 1460 810 1469
rect 162 1426 810 1460
rect 162 1417 810 1426
rect 900 1374 1548 1383
rect 900 1340 1548 1374
rect 900 1331 1548 1340
rect 162 1288 810 1297
rect 162 1254 810 1288
rect 162 1245 810 1254
rect 900 1202 1548 1211
rect 900 1168 1548 1202
rect 900 1159 1548 1168
rect 162 1116 810 1125
rect 162 1082 810 1116
rect 162 1073 810 1082
rect 900 1030 1548 1039
rect 900 996 1548 1030
rect 900 987 1548 996
rect 162 944 810 953
rect 162 910 810 944
rect 162 901 810 910
rect 900 858 1548 867
rect 900 824 1548 858
rect 900 815 1548 824
rect 162 772 810 781
rect 162 738 810 772
rect 162 729 810 738
rect 900 686 1548 695
rect 900 652 1548 686
rect 900 643 1548 652
rect 162 600 810 609
rect 162 566 810 600
rect 162 557 810 566
rect 900 514 1548 523
rect 900 480 1548 514
rect 900 471 1548 480
rect 162 428 810 437
rect 162 394 810 428
rect 162 385 810 394
rect 900 342 1548 351
rect 900 308 1548 342
rect 900 299 1548 308
rect 162 256 810 265
rect 162 222 810 256
rect 162 213 810 222
rect 1618 179 1628 21111
rect 1628 179 1662 21111
rect 1662 179 1672 21111
rect 900 170 1548 179
rect 900 136 1548 170
rect 1618 169 1672 179
rect 900 127 1548 136
<< metal2 >>
rect 156 21077 816 21163
rect 156 21025 162 21077
rect 810 21025 816 21077
rect 156 20905 816 21025
rect 156 20853 162 20905
rect 810 20853 816 20905
rect 156 20733 816 20853
rect 156 20681 162 20733
rect 810 20681 816 20733
rect 156 20561 816 20681
rect 156 20509 162 20561
rect 810 20509 816 20561
rect 156 20389 816 20509
rect 156 20337 162 20389
rect 810 20337 816 20389
rect 156 20217 816 20337
rect 156 20165 162 20217
rect 810 20165 816 20217
rect 156 20045 816 20165
rect 156 19993 162 20045
rect 810 19993 816 20045
rect 156 19873 816 19993
rect 156 19821 162 19873
rect 810 19821 816 19873
rect 156 19701 816 19821
rect 156 19649 162 19701
rect 810 19649 816 19701
rect 156 19529 816 19649
rect 156 19477 162 19529
rect 810 19477 816 19529
rect 156 19357 816 19477
rect 156 19305 162 19357
rect 810 19305 816 19357
rect 156 19185 816 19305
rect 156 19133 162 19185
rect 810 19133 816 19185
rect 156 19013 816 19133
rect 156 18961 162 19013
rect 810 18961 816 19013
rect 156 18841 816 18961
rect 156 18789 162 18841
rect 810 18789 816 18841
rect 156 18669 816 18789
rect 156 18617 162 18669
rect 810 18617 816 18669
rect 156 18497 816 18617
rect 156 18445 162 18497
rect 810 18445 816 18497
rect 156 18325 816 18445
rect 156 18273 162 18325
rect 810 18273 816 18325
rect 156 18153 816 18273
rect 156 18101 162 18153
rect 810 18101 816 18153
rect 156 17981 816 18101
rect 156 17929 162 17981
rect 810 17929 816 17981
rect 156 17809 816 17929
rect 156 17757 162 17809
rect 810 17757 816 17809
rect 156 17637 816 17757
rect 156 17585 162 17637
rect 810 17585 816 17637
rect 156 17465 816 17585
rect 156 17413 162 17465
rect 810 17413 816 17465
rect 156 17293 816 17413
rect 156 17241 162 17293
rect 810 17241 816 17293
rect 156 17121 816 17241
rect 156 17069 162 17121
rect 810 17069 816 17121
rect 156 16949 816 17069
rect 156 16897 162 16949
rect 810 16897 816 16949
rect 156 16777 816 16897
rect 156 16725 162 16777
rect 810 16725 816 16777
rect 156 16605 816 16725
rect 156 16553 162 16605
rect 810 16553 816 16605
rect 156 16433 816 16553
rect 156 16381 162 16433
rect 810 16381 816 16433
rect 156 16261 816 16381
rect 156 16209 162 16261
rect 810 16209 816 16261
rect 156 16089 816 16209
rect 156 16037 162 16089
rect 810 16037 816 16089
rect 156 15917 816 16037
rect 156 15865 162 15917
rect 810 15865 816 15917
rect 156 15745 816 15865
rect 156 15693 162 15745
rect 810 15693 816 15745
rect 156 15573 816 15693
rect 156 15521 162 15573
rect 810 15521 816 15573
rect 156 15401 816 15521
rect 156 15349 162 15401
rect 810 15349 816 15401
rect 156 15229 816 15349
rect 156 15177 162 15229
rect 810 15177 816 15229
rect 156 15057 816 15177
rect 156 15005 162 15057
rect 810 15005 816 15057
rect 156 14885 816 15005
rect 156 14833 162 14885
rect 810 14833 816 14885
rect 156 14713 816 14833
rect 156 14661 162 14713
rect 810 14661 816 14713
rect 156 14541 816 14661
rect 156 14489 162 14541
rect 810 14489 816 14541
rect 156 14369 816 14489
rect 156 14317 162 14369
rect 810 14317 816 14369
rect 156 14197 816 14317
rect 156 14145 162 14197
rect 810 14145 816 14197
rect 156 14025 816 14145
rect 156 13973 162 14025
rect 810 13973 816 14025
rect 156 13853 816 13973
rect 156 13801 162 13853
rect 810 13801 816 13853
rect 156 13681 816 13801
rect 156 13629 162 13681
rect 810 13629 816 13681
rect 156 13509 816 13629
rect 156 13457 162 13509
rect 810 13457 816 13509
rect 156 13337 816 13457
rect 156 13285 162 13337
rect 810 13285 816 13337
rect 156 13165 816 13285
rect 156 13113 162 13165
rect 810 13113 816 13165
rect 156 12993 816 13113
rect 156 12941 162 12993
rect 810 12941 816 12993
rect 156 12821 816 12941
rect 156 12769 162 12821
rect 810 12769 816 12821
rect 156 12649 816 12769
rect 156 12597 162 12649
rect 810 12597 816 12649
rect 156 12477 816 12597
rect 156 12425 162 12477
rect 810 12425 816 12477
rect 156 12305 816 12425
rect 156 12253 162 12305
rect 810 12253 816 12305
rect 156 12133 816 12253
rect 156 12081 162 12133
rect 810 12081 816 12133
rect 156 11961 816 12081
rect 156 11909 162 11961
rect 810 11909 816 11961
rect 156 11789 816 11909
rect 156 11737 162 11789
rect 810 11737 816 11789
rect 156 11617 816 11737
rect 156 11565 162 11617
rect 810 11565 816 11617
rect 156 11445 816 11565
rect 156 11393 162 11445
rect 810 11393 816 11445
rect 156 11273 816 11393
rect 156 11221 162 11273
rect 810 11221 816 11273
rect 156 11101 816 11221
rect 156 11049 162 11101
rect 810 11049 816 11101
rect 156 10929 816 11049
rect 156 10877 162 10929
rect 810 10877 816 10929
rect 156 10757 816 10877
rect 156 10705 162 10757
rect 810 10705 816 10757
rect 156 10585 816 10705
rect 156 10533 162 10585
rect 810 10533 816 10585
rect 156 10413 816 10533
rect 156 10361 162 10413
rect 810 10361 816 10413
rect 156 10241 816 10361
rect 156 10189 162 10241
rect 810 10189 816 10241
rect 156 10069 816 10189
rect 156 10017 162 10069
rect 810 10017 816 10069
rect 156 9897 816 10017
rect 156 9845 162 9897
rect 810 9845 816 9897
rect 156 9725 816 9845
rect 156 9673 162 9725
rect 810 9673 816 9725
rect 156 9553 816 9673
rect 156 9501 162 9553
rect 810 9501 816 9553
rect 156 9381 816 9501
rect 156 9329 162 9381
rect 810 9329 816 9381
rect 156 9209 816 9329
rect 156 9157 162 9209
rect 810 9157 816 9209
rect 156 9037 816 9157
rect 156 8985 162 9037
rect 810 8985 816 9037
rect 156 8865 816 8985
rect 156 8813 162 8865
rect 810 8813 816 8865
rect 156 8693 816 8813
rect 156 8641 162 8693
rect 810 8641 816 8693
rect 156 8521 816 8641
rect 156 8469 162 8521
rect 810 8469 816 8521
rect 156 8349 816 8469
rect 156 8297 162 8349
rect 810 8297 816 8349
rect 156 8177 816 8297
rect 156 8125 162 8177
rect 810 8125 816 8177
rect 156 8005 816 8125
rect 156 7953 162 8005
rect 810 7953 816 8005
rect 156 7833 816 7953
rect 156 7781 162 7833
rect 810 7781 816 7833
rect 156 7661 816 7781
rect 156 7609 162 7661
rect 810 7609 816 7661
rect 156 7489 816 7609
rect 156 7437 162 7489
rect 810 7437 816 7489
rect 156 7317 816 7437
rect 156 7265 162 7317
rect 810 7265 816 7317
rect 156 7145 816 7265
rect 156 7093 162 7145
rect 810 7093 816 7145
rect 156 6973 816 7093
rect 156 6921 162 6973
rect 810 6921 816 6973
rect 156 6801 816 6921
rect 156 6749 162 6801
rect 810 6749 816 6801
rect 156 6629 816 6749
rect 156 6577 162 6629
rect 810 6577 816 6629
rect 156 6457 816 6577
rect 156 6405 162 6457
rect 810 6405 816 6457
rect 156 6285 816 6405
rect 156 6233 162 6285
rect 810 6233 816 6285
rect 156 6113 816 6233
rect 156 6061 162 6113
rect 810 6061 816 6113
rect 156 5941 816 6061
rect 156 5889 162 5941
rect 810 5889 816 5941
rect 156 5769 816 5889
rect 156 5717 162 5769
rect 810 5717 816 5769
rect 156 5597 816 5717
rect 156 5545 162 5597
rect 810 5545 816 5597
rect 156 5425 816 5545
rect 156 5373 162 5425
rect 810 5373 816 5425
rect 156 5253 816 5373
rect 156 5201 162 5253
rect 810 5201 816 5253
rect 156 5081 816 5201
rect 156 5029 162 5081
rect 810 5029 816 5081
rect 156 4909 816 5029
rect 156 4857 162 4909
rect 810 4857 816 4909
rect 156 4737 816 4857
rect 156 4685 162 4737
rect 810 4685 816 4737
rect 156 4565 816 4685
rect 156 4513 162 4565
rect 810 4513 816 4565
rect 156 4393 816 4513
rect 156 4341 162 4393
rect 810 4341 816 4393
rect 156 4221 816 4341
rect 156 4169 162 4221
rect 810 4169 816 4221
rect 156 4049 816 4169
rect 156 3997 162 4049
rect 810 3997 816 4049
rect 156 3877 816 3997
rect 156 3825 162 3877
rect 810 3825 816 3877
rect 156 3705 816 3825
rect 156 3653 162 3705
rect 810 3653 816 3705
rect 156 3533 816 3653
rect 156 3481 162 3533
rect 810 3481 816 3533
rect 156 3361 816 3481
rect 156 3309 162 3361
rect 810 3309 816 3361
rect 156 3189 816 3309
rect 156 3137 162 3189
rect 810 3137 816 3189
rect 156 3017 816 3137
rect 156 2965 162 3017
rect 810 2965 816 3017
rect 156 2845 816 2965
rect 156 2793 162 2845
rect 810 2793 816 2845
rect 156 2673 816 2793
rect 156 2621 162 2673
rect 810 2621 816 2673
rect 156 2501 816 2621
rect 156 2449 162 2501
rect 810 2449 816 2501
rect 156 2329 816 2449
rect 156 2277 162 2329
rect 810 2277 816 2329
rect 156 2157 816 2277
rect 156 2105 162 2157
rect 810 2105 816 2157
rect 156 1985 816 2105
rect 156 1933 162 1985
rect 810 1933 816 1985
rect 156 1813 816 1933
rect 156 1761 162 1813
rect 810 1761 816 1813
rect 156 1641 816 1761
rect 156 1589 162 1641
rect 810 1589 816 1641
rect 156 1469 816 1589
rect 156 1417 162 1469
rect 810 1417 816 1469
rect 156 1297 816 1417
rect 156 1245 162 1297
rect 810 1245 816 1297
rect 156 1125 816 1245
rect 156 1073 162 1125
rect 810 1073 816 1125
rect 156 953 816 1073
rect 156 901 162 953
rect 810 901 816 953
rect 156 781 816 901
rect 156 729 162 781
rect 810 729 816 781
rect 156 609 816 729
rect 156 557 162 609
rect 810 557 816 609
rect 156 437 816 557
rect 156 385 162 437
rect 810 385 816 437
rect 156 265 816 385
rect 156 213 162 265
rect 810 213 816 265
rect 156 127 816 213
rect 894 21111 900 21163
rect 1548 21111 1554 21163
rect 894 20991 1554 21111
rect 894 20939 900 20991
rect 1548 20939 1554 20991
rect 894 20819 1554 20939
rect 894 20767 900 20819
rect 1548 20767 1554 20819
rect 894 20647 1554 20767
rect 894 20595 900 20647
rect 1548 20595 1554 20647
rect 894 20475 1554 20595
rect 894 20423 900 20475
rect 1548 20423 1554 20475
rect 894 20303 1554 20423
rect 894 20251 900 20303
rect 1548 20251 1554 20303
rect 894 20131 1554 20251
rect 894 20079 900 20131
rect 1548 20079 1554 20131
rect 894 19959 1554 20079
rect 894 19907 900 19959
rect 1548 19907 1554 19959
rect 894 19787 1554 19907
rect 894 19735 900 19787
rect 1548 19735 1554 19787
rect 894 19615 1554 19735
rect 894 19563 900 19615
rect 1548 19563 1554 19615
rect 894 19443 1554 19563
rect 894 19391 900 19443
rect 1548 19391 1554 19443
rect 894 19271 1554 19391
rect 894 19219 900 19271
rect 1548 19219 1554 19271
rect 894 19099 1554 19219
rect 894 19047 900 19099
rect 1548 19047 1554 19099
rect 894 18927 1554 19047
rect 894 18875 900 18927
rect 1548 18875 1554 18927
rect 894 18755 1554 18875
rect 894 18703 900 18755
rect 1548 18703 1554 18755
rect 894 18583 1554 18703
rect 894 18531 900 18583
rect 1548 18531 1554 18583
rect 894 18411 1554 18531
rect 894 18359 900 18411
rect 1548 18359 1554 18411
rect 894 18239 1554 18359
rect 894 18187 900 18239
rect 1548 18187 1554 18239
rect 894 18067 1554 18187
rect 894 18015 900 18067
rect 1548 18015 1554 18067
rect 894 17895 1554 18015
rect 894 17843 900 17895
rect 1548 17843 1554 17895
rect 894 17723 1554 17843
rect 894 17671 900 17723
rect 1548 17671 1554 17723
rect 894 17551 1554 17671
rect 894 17499 900 17551
rect 1548 17499 1554 17551
rect 894 17379 1554 17499
rect 894 17327 900 17379
rect 1548 17327 1554 17379
rect 894 17207 1554 17327
rect 894 17155 900 17207
rect 1548 17155 1554 17207
rect 894 17035 1554 17155
rect 894 16983 900 17035
rect 1548 16983 1554 17035
rect 894 16863 1554 16983
rect 894 16811 900 16863
rect 1548 16811 1554 16863
rect 894 16691 1554 16811
rect 894 16639 900 16691
rect 1548 16639 1554 16691
rect 894 16519 1554 16639
rect 894 16467 900 16519
rect 1548 16467 1554 16519
rect 894 16347 1554 16467
rect 894 16295 900 16347
rect 1548 16295 1554 16347
rect 894 16175 1554 16295
rect 894 16123 900 16175
rect 1548 16123 1554 16175
rect 894 16003 1554 16123
rect 894 15951 900 16003
rect 1548 15951 1554 16003
rect 894 15831 1554 15951
rect 894 15779 900 15831
rect 1548 15779 1554 15831
rect 894 15659 1554 15779
rect 894 15607 900 15659
rect 1548 15607 1554 15659
rect 894 15487 1554 15607
rect 894 15435 900 15487
rect 1548 15435 1554 15487
rect 894 15315 1554 15435
rect 894 15263 900 15315
rect 1548 15263 1554 15315
rect 894 15143 1554 15263
rect 894 15091 900 15143
rect 1548 15091 1554 15143
rect 894 14971 1554 15091
rect 894 14919 900 14971
rect 1548 14919 1554 14971
rect 894 14799 1554 14919
rect 894 14747 900 14799
rect 1548 14747 1554 14799
rect 894 14627 1554 14747
rect 894 14575 900 14627
rect 1548 14575 1554 14627
rect 894 14455 1554 14575
rect 894 14403 900 14455
rect 1548 14403 1554 14455
rect 894 14283 1554 14403
rect 894 14231 900 14283
rect 1548 14231 1554 14283
rect 894 14111 1554 14231
rect 894 14059 900 14111
rect 1548 14059 1554 14111
rect 894 13939 1554 14059
rect 894 13887 900 13939
rect 1548 13887 1554 13939
rect 894 13767 1554 13887
rect 894 13715 900 13767
rect 1548 13715 1554 13767
rect 894 13595 1554 13715
rect 894 13543 900 13595
rect 1548 13543 1554 13595
rect 894 13423 1554 13543
rect 894 13371 900 13423
rect 1548 13371 1554 13423
rect 894 13251 1554 13371
rect 894 13199 900 13251
rect 1548 13199 1554 13251
rect 894 13079 1554 13199
rect 894 13027 900 13079
rect 1548 13027 1554 13079
rect 894 12907 1554 13027
rect 894 12855 900 12907
rect 1548 12855 1554 12907
rect 894 12735 1554 12855
rect 894 12683 900 12735
rect 1548 12683 1554 12735
rect 894 12563 1554 12683
rect 894 12511 900 12563
rect 1548 12511 1554 12563
rect 894 12391 1554 12511
rect 894 12339 900 12391
rect 1548 12339 1554 12391
rect 894 12219 1554 12339
rect 894 12167 900 12219
rect 1548 12167 1554 12219
rect 894 12047 1554 12167
rect 894 11995 900 12047
rect 1548 11995 1554 12047
rect 894 11875 1554 11995
rect 894 11823 900 11875
rect 1548 11823 1554 11875
rect 894 11703 1554 11823
rect 894 11651 900 11703
rect 1548 11651 1554 11703
rect 894 11531 1554 11651
rect 894 11479 900 11531
rect 1548 11479 1554 11531
rect 894 11359 1554 11479
rect 894 11307 900 11359
rect 1548 11307 1554 11359
rect 894 11187 1554 11307
rect 894 11135 900 11187
rect 1548 11135 1554 11187
rect 894 11015 1554 11135
rect 894 10963 900 11015
rect 1548 10963 1554 11015
rect 894 10843 1554 10963
rect 894 10791 900 10843
rect 1548 10791 1554 10843
rect 894 10671 1554 10791
rect 894 10619 900 10671
rect 1548 10619 1554 10671
rect 894 10499 1554 10619
rect 894 10447 900 10499
rect 1548 10447 1554 10499
rect 894 10327 1554 10447
rect 894 10275 900 10327
rect 1548 10275 1554 10327
rect 894 10155 1554 10275
rect 894 10103 900 10155
rect 1548 10103 1554 10155
rect 894 9983 1554 10103
rect 894 9931 900 9983
rect 1548 9931 1554 9983
rect 894 9811 1554 9931
rect 894 9759 900 9811
rect 1548 9759 1554 9811
rect 894 9639 1554 9759
rect 894 9587 900 9639
rect 1548 9587 1554 9639
rect 894 9467 1554 9587
rect 894 9415 900 9467
rect 1548 9415 1554 9467
rect 894 9295 1554 9415
rect 894 9243 900 9295
rect 1548 9243 1554 9295
rect 894 9123 1554 9243
rect 894 9071 900 9123
rect 1548 9071 1554 9123
rect 894 8951 1554 9071
rect 894 8899 900 8951
rect 1548 8899 1554 8951
rect 894 8779 1554 8899
rect 894 8727 900 8779
rect 1548 8727 1554 8779
rect 894 8607 1554 8727
rect 894 8555 900 8607
rect 1548 8555 1554 8607
rect 894 8435 1554 8555
rect 894 8383 900 8435
rect 1548 8383 1554 8435
rect 894 8263 1554 8383
rect 894 8211 900 8263
rect 1548 8211 1554 8263
rect 894 8091 1554 8211
rect 894 8039 900 8091
rect 1548 8039 1554 8091
rect 894 7919 1554 8039
rect 894 7867 900 7919
rect 1548 7867 1554 7919
rect 894 7747 1554 7867
rect 894 7695 900 7747
rect 1548 7695 1554 7747
rect 894 7575 1554 7695
rect 894 7523 900 7575
rect 1548 7523 1554 7575
rect 894 7403 1554 7523
rect 894 7351 900 7403
rect 1548 7351 1554 7403
rect 894 7231 1554 7351
rect 894 7179 900 7231
rect 1548 7179 1554 7231
rect 894 7059 1554 7179
rect 894 7007 900 7059
rect 1548 7007 1554 7059
rect 894 6887 1554 7007
rect 894 6835 900 6887
rect 1548 6835 1554 6887
rect 894 6715 1554 6835
rect 894 6663 900 6715
rect 1548 6663 1554 6715
rect 894 6543 1554 6663
rect 894 6491 900 6543
rect 1548 6491 1554 6543
rect 894 6371 1554 6491
rect 894 6319 900 6371
rect 1548 6319 1554 6371
rect 894 6199 1554 6319
rect 894 6147 900 6199
rect 1548 6147 1554 6199
rect 894 6027 1554 6147
rect 894 5975 900 6027
rect 1548 5975 1554 6027
rect 894 5855 1554 5975
rect 894 5803 900 5855
rect 1548 5803 1554 5855
rect 894 5683 1554 5803
rect 894 5631 900 5683
rect 1548 5631 1554 5683
rect 894 5511 1554 5631
rect 894 5459 900 5511
rect 1548 5459 1554 5511
rect 894 5339 1554 5459
rect 894 5287 900 5339
rect 1548 5287 1554 5339
rect 894 5167 1554 5287
rect 894 5115 900 5167
rect 1548 5115 1554 5167
rect 894 4995 1554 5115
rect 894 4943 900 4995
rect 1548 4943 1554 4995
rect 894 4823 1554 4943
rect 894 4771 900 4823
rect 1548 4771 1554 4823
rect 894 4651 1554 4771
rect 894 4599 900 4651
rect 1548 4599 1554 4651
rect 894 4479 1554 4599
rect 894 4427 900 4479
rect 1548 4427 1554 4479
rect 894 4307 1554 4427
rect 894 4255 900 4307
rect 1548 4255 1554 4307
rect 894 4135 1554 4255
rect 894 4083 900 4135
rect 1548 4083 1554 4135
rect 894 3963 1554 4083
rect 894 3911 900 3963
rect 1548 3911 1554 3963
rect 894 3791 1554 3911
rect 894 3739 900 3791
rect 1548 3739 1554 3791
rect 894 3619 1554 3739
rect 894 3567 900 3619
rect 1548 3567 1554 3619
rect 894 3447 1554 3567
rect 894 3395 900 3447
rect 1548 3395 1554 3447
rect 894 3275 1554 3395
rect 894 3223 900 3275
rect 1548 3223 1554 3275
rect 894 3103 1554 3223
rect 894 3051 900 3103
rect 1548 3051 1554 3103
rect 894 2931 1554 3051
rect 894 2879 900 2931
rect 1548 2879 1554 2931
rect 894 2759 1554 2879
rect 894 2707 900 2759
rect 1548 2707 1554 2759
rect 894 2587 1554 2707
rect 894 2535 900 2587
rect 1548 2535 1554 2587
rect 894 2415 1554 2535
rect 894 2363 900 2415
rect 1548 2363 1554 2415
rect 894 2243 1554 2363
rect 894 2191 900 2243
rect 1548 2191 1554 2243
rect 894 2071 1554 2191
rect 894 2019 900 2071
rect 1548 2019 1554 2071
rect 894 1899 1554 2019
rect 894 1847 900 1899
rect 1548 1847 1554 1899
rect 894 1727 1554 1847
rect 894 1675 900 1727
rect 1548 1675 1554 1727
rect 894 1555 1554 1675
rect 894 1503 900 1555
rect 1548 1503 1554 1555
rect 894 1383 1554 1503
rect 894 1331 900 1383
rect 1548 1331 1554 1383
rect 894 1211 1554 1331
rect 894 1159 900 1211
rect 1548 1159 1554 1211
rect 894 1039 1554 1159
rect 894 987 900 1039
rect 1548 987 1554 1039
rect 894 867 1554 987
rect 894 815 900 867
rect 1548 815 1554 867
rect 894 695 1554 815
rect 894 643 900 695
rect 1548 643 1554 695
rect 894 523 1554 643
rect 894 471 900 523
rect 1548 471 1554 523
rect 894 351 1554 471
rect 894 299 900 351
rect 1548 299 1554 351
rect 894 179 1554 299
rect 894 127 900 179
rect 1548 127 1554 179
rect 1618 21121 1672 21127
rect 1618 163 1672 169
<< end >>
