magic
tech sky130A
magscale 1 2
timestamp 1712480545
<< error_p >>
rect -1311 531 -1249 537
rect -1183 531 -1121 537
rect -1055 531 -993 537
rect -927 531 -865 537
rect -799 531 -737 537
rect -671 531 -609 537
rect -543 531 -481 537
rect -415 531 -353 537
rect -287 531 -225 537
rect -159 531 -97 537
rect -31 531 31 537
rect 97 531 159 537
rect 225 531 287 537
rect 353 531 415 537
rect 481 531 543 537
rect 609 531 671 537
rect 737 531 799 537
rect 865 531 927 537
rect 993 531 1055 537
rect 1121 531 1183 537
rect 1249 531 1311 537
rect -1311 497 -1299 531
rect -1183 497 -1171 531
rect -1055 497 -1043 531
rect -927 497 -915 531
rect -799 497 -787 531
rect -671 497 -659 531
rect -543 497 -531 531
rect -415 497 -403 531
rect -287 497 -275 531
rect -159 497 -147 531
rect -31 497 -19 531
rect 97 497 109 531
rect 225 497 237 531
rect 353 497 365 531
rect 481 497 493 531
rect 609 497 621 531
rect 737 497 749 531
rect 865 497 877 531
rect 993 497 1005 531
rect 1121 497 1133 531
rect 1249 497 1261 531
rect -1311 491 -1249 497
rect -1183 491 -1121 497
rect -1055 491 -993 497
rect -927 491 -865 497
rect -799 491 -737 497
rect -671 491 -609 497
rect -543 491 -481 497
rect -415 491 -353 497
rect -287 491 -225 497
rect -159 491 -97 497
rect -31 491 31 497
rect 97 491 159 497
rect 225 491 287 497
rect 353 491 415 497
rect 481 491 543 497
rect 609 491 671 497
rect 737 491 799 497
rect 865 491 927 497
rect 993 491 1055 497
rect 1121 491 1183 497
rect 1249 491 1311 497
rect -1311 -497 -1249 -491
rect -1183 -497 -1121 -491
rect -1055 -497 -993 -491
rect -927 -497 -865 -491
rect -799 -497 -737 -491
rect -671 -497 -609 -491
rect -543 -497 -481 -491
rect -415 -497 -353 -491
rect -287 -497 -225 -491
rect -159 -497 -97 -491
rect -31 -497 31 -491
rect 97 -497 159 -491
rect 225 -497 287 -491
rect 353 -497 415 -491
rect 481 -497 543 -491
rect 609 -497 671 -491
rect 737 -497 799 -491
rect 865 -497 927 -491
rect 993 -497 1055 -491
rect 1121 -497 1183 -491
rect 1249 -497 1311 -491
rect -1311 -531 -1299 -497
rect -1183 -531 -1171 -497
rect -1055 -531 -1043 -497
rect -927 -531 -915 -497
rect -799 -531 -787 -497
rect -671 -531 -659 -497
rect -543 -531 -531 -497
rect -415 -531 -403 -497
rect -287 -531 -275 -497
rect -159 -531 -147 -497
rect -31 -531 -19 -497
rect 97 -531 109 -497
rect 225 -531 237 -497
rect 353 -531 365 -497
rect 481 -531 493 -497
rect 609 -531 621 -497
rect 737 -531 749 -497
rect 865 -531 877 -497
rect 993 -531 1005 -497
rect 1121 -531 1133 -497
rect 1249 -531 1261 -497
rect -1311 -537 -1249 -531
rect -1183 -537 -1121 -531
rect -1055 -537 -993 -531
rect -927 -537 -865 -531
rect -799 -537 -737 -531
rect -671 -537 -609 -531
rect -543 -537 -481 -531
rect -415 -537 -353 -531
rect -287 -537 -225 -531
rect -159 -537 -97 -531
rect -31 -537 31 -531
rect 97 -537 159 -531
rect 225 -537 287 -531
rect 353 -537 415 -531
rect 481 -537 543 -531
rect 609 -537 671 -531
rect 737 -537 799 -531
rect 865 -537 927 -531
rect 993 -537 1055 -531
rect 1121 -537 1183 -531
rect 1249 -537 1311 -531
<< nwell >>
rect -1511 -669 1511 669
<< pmoslvt >>
rect -1315 -450 -1245 450
rect -1187 -450 -1117 450
rect -1059 -450 -989 450
rect -931 -450 -861 450
rect -803 -450 -733 450
rect -675 -450 -605 450
rect -547 -450 -477 450
rect -419 -450 -349 450
rect -291 -450 -221 450
rect -163 -450 -93 450
rect -35 -450 35 450
rect 93 -450 163 450
rect 221 -450 291 450
rect 349 -450 419 450
rect 477 -450 547 450
rect 605 -450 675 450
rect 733 -450 803 450
rect 861 -450 931 450
rect 989 -450 1059 450
rect 1117 -450 1187 450
rect 1245 -450 1315 450
<< pdiff >>
rect -1373 438 -1315 450
rect -1373 -438 -1361 438
rect -1327 -438 -1315 438
rect -1373 -450 -1315 -438
rect -1245 438 -1187 450
rect -1245 -438 -1233 438
rect -1199 -438 -1187 438
rect -1245 -450 -1187 -438
rect -1117 438 -1059 450
rect -1117 -438 -1105 438
rect -1071 -438 -1059 438
rect -1117 -450 -1059 -438
rect -989 438 -931 450
rect -989 -438 -977 438
rect -943 -438 -931 438
rect -989 -450 -931 -438
rect -861 438 -803 450
rect -861 -438 -849 438
rect -815 -438 -803 438
rect -861 -450 -803 -438
rect -733 438 -675 450
rect -733 -438 -721 438
rect -687 -438 -675 438
rect -733 -450 -675 -438
rect -605 438 -547 450
rect -605 -438 -593 438
rect -559 -438 -547 438
rect -605 -450 -547 -438
rect -477 438 -419 450
rect -477 -438 -465 438
rect -431 -438 -419 438
rect -477 -450 -419 -438
rect -349 438 -291 450
rect -349 -438 -337 438
rect -303 -438 -291 438
rect -349 -450 -291 -438
rect -221 438 -163 450
rect -221 -438 -209 438
rect -175 -438 -163 438
rect -221 -450 -163 -438
rect -93 438 -35 450
rect -93 -438 -81 438
rect -47 -438 -35 438
rect -93 -450 -35 -438
rect 35 438 93 450
rect 35 -438 47 438
rect 81 -438 93 438
rect 35 -450 93 -438
rect 163 438 221 450
rect 163 -438 175 438
rect 209 -438 221 438
rect 163 -450 221 -438
rect 291 438 349 450
rect 291 -438 303 438
rect 337 -438 349 438
rect 291 -450 349 -438
rect 419 438 477 450
rect 419 -438 431 438
rect 465 -438 477 438
rect 419 -450 477 -438
rect 547 438 605 450
rect 547 -438 559 438
rect 593 -438 605 438
rect 547 -450 605 -438
rect 675 438 733 450
rect 675 -438 687 438
rect 721 -438 733 438
rect 675 -450 733 -438
rect 803 438 861 450
rect 803 -438 815 438
rect 849 -438 861 438
rect 803 -450 861 -438
rect 931 438 989 450
rect 931 -438 943 438
rect 977 -438 989 438
rect 931 -450 989 -438
rect 1059 438 1117 450
rect 1059 -438 1071 438
rect 1105 -438 1117 438
rect 1059 -450 1117 -438
rect 1187 438 1245 450
rect 1187 -438 1199 438
rect 1233 -438 1245 438
rect 1187 -450 1245 -438
rect 1315 438 1373 450
rect 1315 -438 1327 438
rect 1361 -438 1373 438
rect 1315 -450 1373 -438
<< pdiffc >>
rect -1361 -438 -1327 438
rect -1233 -438 -1199 438
rect -1105 -438 -1071 438
rect -977 -438 -943 438
rect -849 -438 -815 438
rect -721 -438 -687 438
rect -593 -438 -559 438
rect -465 -438 -431 438
rect -337 -438 -303 438
rect -209 -438 -175 438
rect -81 -438 -47 438
rect 47 -438 81 438
rect 175 -438 209 438
rect 303 -438 337 438
rect 431 -438 465 438
rect 559 -438 593 438
rect 687 -438 721 438
rect 815 -438 849 438
rect 943 -438 977 438
rect 1071 -438 1105 438
rect 1199 -438 1233 438
rect 1327 -438 1361 438
<< nsubdiff >>
rect -1475 599 -1379 633
rect 1379 599 1475 633
rect -1475 537 -1441 599
rect 1441 537 1475 599
rect -1475 -599 -1441 -537
rect 1441 -599 1475 -537
rect -1475 -633 -1379 -599
rect 1379 -633 1475 -599
<< nsubdiffcont >>
rect -1379 599 1379 633
rect -1475 -537 -1441 537
rect 1441 -537 1475 537
rect -1379 -633 1379 -599
<< poly >>
rect -1315 531 -1245 547
rect -1315 497 -1299 531
rect -1261 497 -1245 531
rect -1315 450 -1245 497
rect -1187 531 -1117 547
rect -1187 497 -1171 531
rect -1133 497 -1117 531
rect -1187 450 -1117 497
rect -1059 531 -989 547
rect -1059 497 -1043 531
rect -1005 497 -989 531
rect -1059 450 -989 497
rect -931 531 -861 547
rect -931 497 -915 531
rect -877 497 -861 531
rect -931 450 -861 497
rect -803 531 -733 547
rect -803 497 -787 531
rect -749 497 -733 531
rect -803 450 -733 497
rect -675 531 -605 547
rect -675 497 -659 531
rect -621 497 -605 531
rect -675 450 -605 497
rect -547 531 -477 547
rect -547 497 -531 531
rect -493 497 -477 531
rect -547 450 -477 497
rect -419 531 -349 547
rect -419 497 -403 531
rect -365 497 -349 531
rect -419 450 -349 497
rect -291 531 -221 547
rect -291 497 -275 531
rect -237 497 -221 531
rect -291 450 -221 497
rect -163 531 -93 547
rect -163 497 -147 531
rect -109 497 -93 531
rect -163 450 -93 497
rect -35 531 35 547
rect -35 497 -19 531
rect 19 497 35 531
rect -35 450 35 497
rect 93 531 163 547
rect 93 497 109 531
rect 147 497 163 531
rect 93 450 163 497
rect 221 531 291 547
rect 221 497 237 531
rect 275 497 291 531
rect 221 450 291 497
rect 349 531 419 547
rect 349 497 365 531
rect 403 497 419 531
rect 349 450 419 497
rect 477 531 547 547
rect 477 497 493 531
rect 531 497 547 531
rect 477 450 547 497
rect 605 531 675 547
rect 605 497 621 531
rect 659 497 675 531
rect 605 450 675 497
rect 733 531 803 547
rect 733 497 749 531
rect 787 497 803 531
rect 733 450 803 497
rect 861 531 931 547
rect 861 497 877 531
rect 915 497 931 531
rect 861 450 931 497
rect 989 531 1059 547
rect 989 497 1005 531
rect 1043 497 1059 531
rect 989 450 1059 497
rect 1117 531 1187 547
rect 1117 497 1133 531
rect 1171 497 1187 531
rect 1117 450 1187 497
rect 1245 531 1315 547
rect 1245 497 1261 531
rect 1299 497 1315 531
rect 1245 450 1315 497
rect -1315 -497 -1245 -450
rect -1315 -531 -1299 -497
rect -1261 -531 -1245 -497
rect -1315 -547 -1245 -531
rect -1187 -497 -1117 -450
rect -1187 -531 -1171 -497
rect -1133 -531 -1117 -497
rect -1187 -547 -1117 -531
rect -1059 -497 -989 -450
rect -1059 -531 -1043 -497
rect -1005 -531 -989 -497
rect -1059 -547 -989 -531
rect -931 -497 -861 -450
rect -931 -531 -915 -497
rect -877 -531 -861 -497
rect -931 -547 -861 -531
rect -803 -497 -733 -450
rect -803 -531 -787 -497
rect -749 -531 -733 -497
rect -803 -547 -733 -531
rect -675 -497 -605 -450
rect -675 -531 -659 -497
rect -621 -531 -605 -497
rect -675 -547 -605 -531
rect -547 -497 -477 -450
rect -547 -531 -531 -497
rect -493 -531 -477 -497
rect -547 -547 -477 -531
rect -419 -497 -349 -450
rect -419 -531 -403 -497
rect -365 -531 -349 -497
rect -419 -547 -349 -531
rect -291 -497 -221 -450
rect -291 -531 -275 -497
rect -237 -531 -221 -497
rect -291 -547 -221 -531
rect -163 -497 -93 -450
rect -163 -531 -147 -497
rect -109 -531 -93 -497
rect -163 -547 -93 -531
rect -35 -497 35 -450
rect -35 -531 -19 -497
rect 19 -531 35 -497
rect -35 -547 35 -531
rect 93 -497 163 -450
rect 93 -531 109 -497
rect 147 -531 163 -497
rect 93 -547 163 -531
rect 221 -497 291 -450
rect 221 -531 237 -497
rect 275 -531 291 -497
rect 221 -547 291 -531
rect 349 -497 419 -450
rect 349 -531 365 -497
rect 403 -531 419 -497
rect 349 -547 419 -531
rect 477 -497 547 -450
rect 477 -531 493 -497
rect 531 -531 547 -497
rect 477 -547 547 -531
rect 605 -497 675 -450
rect 605 -531 621 -497
rect 659 -531 675 -497
rect 605 -547 675 -531
rect 733 -497 803 -450
rect 733 -531 749 -497
rect 787 -531 803 -497
rect 733 -547 803 -531
rect 861 -497 931 -450
rect 861 -531 877 -497
rect 915 -531 931 -497
rect 861 -547 931 -531
rect 989 -497 1059 -450
rect 989 -531 1005 -497
rect 1043 -531 1059 -497
rect 989 -547 1059 -531
rect 1117 -497 1187 -450
rect 1117 -531 1133 -497
rect 1171 -531 1187 -497
rect 1117 -547 1187 -531
rect 1245 -497 1315 -450
rect 1245 -531 1261 -497
rect 1299 -531 1315 -497
rect 1245 -547 1315 -531
<< polycont >>
rect -1299 497 -1261 531
rect -1171 497 -1133 531
rect -1043 497 -1005 531
rect -915 497 -877 531
rect -787 497 -749 531
rect -659 497 -621 531
rect -531 497 -493 531
rect -403 497 -365 531
rect -275 497 -237 531
rect -147 497 -109 531
rect -19 497 19 531
rect 109 497 147 531
rect 237 497 275 531
rect 365 497 403 531
rect 493 497 531 531
rect 621 497 659 531
rect 749 497 787 531
rect 877 497 915 531
rect 1005 497 1043 531
rect 1133 497 1171 531
rect 1261 497 1299 531
rect -1299 -531 -1261 -497
rect -1171 -531 -1133 -497
rect -1043 -531 -1005 -497
rect -915 -531 -877 -497
rect -787 -531 -749 -497
rect -659 -531 -621 -497
rect -531 -531 -493 -497
rect -403 -531 -365 -497
rect -275 -531 -237 -497
rect -147 -531 -109 -497
rect -19 -531 19 -497
rect 109 -531 147 -497
rect 237 -531 275 -497
rect 365 -531 403 -497
rect 493 -531 531 -497
rect 621 -531 659 -497
rect 749 -531 787 -497
rect 877 -531 915 -497
rect 1005 -531 1043 -497
rect 1133 -531 1171 -497
rect 1261 -531 1299 -497
<< locali >>
rect -1475 599 -1379 633
rect 1379 599 1475 633
rect -1475 537 -1441 599
rect 1441 537 1475 599
rect -1315 497 -1299 531
rect -1261 497 -1245 531
rect -1187 497 -1171 531
rect -1133 497 -1117 531
rect -1059 497 -1043 531
rect -1005 497 -989 531
rect -931 497 -915 531
rect -877 497 -861 531
rect -803 497 -787 531
rect -749 497 -733 531
rect -675 497 -659 531
rect -621 497 -605 531
rect -547 497 -531 531
rect -493 497 -477 531
rect -419 497 -403 531
rect -365 497 -349 531
rect -291 497 -275 531
rect -237 497 -221 531
rect -163 497 -147 531
rect -109 497 -93 531
rect -35 497 -19 531
rect 19 497 35 531
rect 93 497 109 531
rect 147 497 163 531
rect 221 497 237 531
rect 275 497 291 531
rect 349 497 365 531
rect 403 497 419 531
rect 477 497 493 531
rect 531 497 547 531
rect 605 497 621 531
rect 659 497 675 531
rect 733 497 749 531
rect 787 497 803 531
rect 861 497 877 531
rect 915 497 931 531
rect 989 497 1005 531
rect 1043 497 1059 531
rect 1117 497 1133 531
rect 1171 497 1187 531
rect 1245 497 1261 531
rect 1299 497 1315 531
rect -1361 438 -1327 454
rect -1361 -454 -1327 -438
rect -1233 438 -1199 454
rect -1233 -454 -1199 -438
rect -1105 438 -1071 454
rect -1105 -454 -1071 -438
rect -977 438 -943 454
rect -977 -454 -943 -438
rect -849 438 -815 454
rect -849 -454 -815 -438
rect -721 438 -687 454
rect -721 -454 -687 -438
rect -593 438 -559 454
rect -593 -454 -559 -438
rect -465 438 -431 454
rect -465 -454 -431 -438
rect -337 438 -303 454
rect -337 -454 -303 -438
rect -209 438 -175 454
rect -209 -454 -175 -438
rect -81 438 -47 454
rect -81 -454 -47 -438
rect 47 438 81 454
rect 47 -454 81 -438
rect 175 438 209 454
rect 175 -454 209 -438
rect 303 438 337 454
rect 303 -454 337 -438
rect 431 438 465 454
rect 431 -454 465 -438
rect 559 438 593 454
rect 559 -454 593 -438
rect 687 438 721 454
rect 687 -454 721 -438
rect 815 438 849 454
rect 815 -454 849 -438
rect 943 438 977 454
rect 943 -454 977 -438
rect 1071 438 1105 454
rect 1071 -454 1105 -438
rect 1199 438 1233 454
rect 1199 -454 1233 -438
rect 1327 438 1361 454
rect 1327 -454 1361 -438
rect -1315 -531 -1299 -497
rect -1261 -531 -1245 -497
rect -1187 -531 -1171 -497
rect -1133 -531 -1117 -497
rect -1059 -531 -1043 -497
rect -1005 -531 -989 -497
rect -931 -531 -915 -497
rect -877 -531 -861 -497
rect -803 -531 -787 -497
rect -749 -531 -733 -497
rect -675 -531 -659 -497
rect -621 -531 -605 -497
rect -547 -531 -531 -497
rect -493 -531 -477 -497
rect -419 -531 -403 -497
rect -365 -531 -349 -497
rect -291 -531 -275 -497
rect -237 -531 -221 -497
rect -163 -531 -147 -497
rect -109 -531 -93 -497
rect -35 -531 -19 -497
rect 19 -531 35 -497
rect 93 -531 109 -497
rect 147 -531 163 -497
rect 221 -531 237 -497
rect 275 -531 291 -497
rect 349 -531 365 -497
rect 403 -531 419 -497
rect 477 -531 493 -497
rect 531 -531 547 -497
rect 605 -531 621 -497
rect 659 -531 675 -497
rect 733 -531 749 -497
rect 787 -531 803 -497
rect 861 -531 877 -497
rect 915 -531 931 -497
rect 989 -531 1005 -497
rect 1043 -531 1059 -497
rect 1117 -531 1133 -497
rect 1171 -531 1187 -497
rect 1245 -531 1261 -497
rect 1299 -531 1315 -497
rect -1475 -599 -1441 -537
rect 1441 -599 1475 -537
rect -1475 -633 -1379 -599
rect 1379 -633 1475 -599
<< viali >>
rect -1299 497 -1261 531
rect -1171 497 -1133 531
rect -1043 497 -1005 531
rect -915 497 -877 531
rect -787 497 -749 531
rect -659 497 -621 531
rect -531 497 -493 531
rect -403 497 -365 531
rect -275 497 -237 531
rect -147 497 -109 531
rect -19 497 19 531
rect 109 497 147 531
rect 237 497 275 531
rect 365 497 403 531
rect 493 497 531 531
rect 621 497 659 531
rect 749 497 787 531
rect 877 497 915 531
rect 1005 497 1043 531
rect 1133 497 1171 531
rect 1261 497 1299 531
rect -1361 -438 -1327 438
rect -1233 -438 -1199 438
rect -1105 -438 -1071 438
rect -977 -438 -943 438
rect -849 -438 -815 438
rect -721 -438 -687 438
rect -593 -438 -559 438
rect -465 -438 -431 438
rect -337 -438 -303 438
rect -209 -438 -175 438
rect -81 -438 -47 438
rect 47 -438 81 438
rect 175 -438 209 438
rect 303 -438 337 438
rect 431 -438 465 438
rect 559 -438 593 438
rect 687 -438 721 438
rect 815 -438 849 438
rect 943 -438 977 438
rect 1071 -438 1105 438
rect 1199 -438 1233 438
rect 1327 -438 1361 438
rect -1299 -531 -1261 -497
rect -1171 -531 -1133 -497
rect -1043 -531 -1005 -497
rect -915 -531 -877 -497
rect -787 -531 -749 -497
rect -659 -531 -621 -497
rect -531 -531 -493 -497
rect -403 -531 -365 -497
rect -275 -531 -237 -497
rect -147 -531 -109 -497
rect -19 -531 19 -497
rect 109 -531 147 -497
rect 237 -531 275 -497
rect 365 -531 403 -497
rect 493 -531 531 -497
rect 621 -531 659 -497
rect 749 -531 787 -497
rect 877 -531 915 -497
rect 1005 -531 1043 -497
rect 1133 -531 1171 -497
rect 1261 -531 1299 -497
<< metal1 >>
rect -1311 531 -1249 537
rect -1311 497 -1299 531
rect -1261 497 -1249 531
rect -1311 491 -1249 497
rect -1183 531 -1121 537
rect -1183 497 -1171 531
rect -1133 497 -1121 531
rect -1183 491 -1121 497
rect -1055 531 -993 537
rect -1055 497 -1043 531
rect -1005 497 -993 531
rect -1055 491 -993 497
rect -927 531 -865 537
rect -927 497 -915 531
rect -877 497 -865 531
rect -927 491 -865 497
rect -799 531 -737 537
rect -799 497 -787 531
rect -749 497 -737 531
rect -799 491 -737 497
rect -671 531 -609 537
rect -671 497 -659 531
rect -621 497 -609 531
rect -671 491 -609 497
rect -543 531 -481 537
rect -543 497 -531 531
rect -493 497 -481 531
rect -543 491 -481 497
rect -415 531 -353 537
rect -415 497 -403 531
rect -365 497 -353 531
rect -415 491 -353 497
rect -287 531 -225 537
rect -287 497 -275 531
rect -237 497 -225 531
rect -287 491 -225 497
rect -159 531 -97 537
rect -159 497 -147 531
rect -109 497 -97 531
rect -159 491 -97 497
rect -31 531 31 537
rect -31 497 -19 531
rect 19 497 31 531
rect -31 491 31 497
rect 97 531 159 537
rect 97 497 109 531
rect 147 497 159 531
rect 97 491 159 497
rect 225 531 287 537
rect 225 497 237 531
rect 275 497 287 531
rect 225 491 287 497
rect 353 531 415 537
rect 353 497 365 531
rect 403 497 415 531
rect 353 491 415 497
rect 481 531 543 537
rect 481 497 493 531
rect 531 497 543 531
rect 481 491 543 497
rect 609 531 671 537
rect 609 497 621 531
rect 659 497 671 531
rect 609 491 671 497
rect 737 531 799 537
rect 737 497 749 531
rect 787 497 799 531
rect 737 491 799 497
rect 865 531 927 537
rect 865 497 877 531
rect 915 497 927 531
rect 865 491 927 497
rect 993 531 1055 537
rect 993 497 1005 531
rect 1043 497 1055 531
rect 993 491 1055 497
rect 1121 531 1183 537
rect 1121 497 1133 531
rect 1171 497 1183 531
rect 1121 491 1183 497
rect 1249 531 1311 537
rect 1249 497 1261 531
rect 1299 497 1311 531
rect 1249 491 1311 497
rect -1367 438 -1321 450
rect -1367 -438 -1361 438
rect -1327 -438 -1321 438
rect -1367 -450 -1321 -438
rect -1239 438 -1193 450
rect -1239 -438 -1233 438
rect -1199 -438 -1193 438
rect -1239 -450 -1193 -438
rect -1111 438 -1065 450
rect -1111 -438 -1105 438
rect -1071 -438 -1065 438
rect -1111 -450 -1065 -438
rect -983 438 -937 450
rect -983 -438 -977 438
rect -943 -438 -937 438
rect -983 -450 -937 -438
rect -855 438 -809 450
rect -855 -438 -849 438
rect -815 -438 -809 438
rect -855 -450 -809 -438
rect -727 438 -681 450
rect -727 -438 -721 438
rect -687 -438 -681 438
rect -727 -450 -681 -438
rect -599 438 -553 450
rect -599 -438 -593 438
rect -559 -438 -553 438
rect -599 -450 -553 -438
rect -471 438 -425 450
rect -471 -438 -465 438
rect -431 -438 -425 438
rect -471 -450 -425 -438
rect -343 438 -297 450
rect -343 -438 -337 438
rect -303 -438 -297 438
rect -343 -450 -297 -438
rect -215 438 -169 450
rect -215 -438 -209 438
rect -175 -438 -169 438
rect -215 -450 -169 -438
rect -87 438 -41 450
rect -87 -438 -81 438
rect -47 -438 -41 438
rect -87 -450 -41 -438
rect 41 438 87 450
rect 41 -438 47 438
rect 81 -438 87 438
rect 41 -450 87 -438
rect 169 438 215 450
rect 169 -438 175 438
rect 209 -438 215 438
rect 169 -450 215 -438
rect 297 438 343 450
rect 297 -438 303 438
rect 337 -438 343 438
rect 297 -450 343 -438
rect 425 438 471 450
rect 425 -438 431 438
rect 465 -438 471 438
rect 425 -450 471 -438
rect 553 438 599 450
rect 553 -438 559 438
rect 593 -438 599 438
rect 553 -450 599 -438
rect 681 438 727 450
rect 681 -438 687 438
rect 721 -438 727 438
rect 681 -450 727 -438
rect 809 438 855 450
rect 809 -438 815 438
rect 849 -438 855 438
rect 809 -450 855 -438
rect 937 438 983 450
rect 937 -438 943 438
rect 977 -438 983 438
rect 937 -450 983 -438
rect 1065 438 1111 450
rect 1065 -438 1071 438
rect 1105 -438 1111 438
rect 1065 -450 1111 -438
rect 1193 438 1239 450
rect 1193 -438 1199 438
rect 1233 -438 1239 438
rect 1193 -450 1239 -438
rect 1321 438 1367 450
rect 1321 -438 1327 438
rect 1361 -438 1367 438
rect 1321 -450 1367 -438
rect -1311 -497 -1249 -491
rect -1311 -531 -1299 -497
rect -1261 -531 -1249 -497
rect -1311 -537 -1249 -531
rect -1183 -497 -1121 -491
rect -1183 -531 -1171 -497
rect -1133 -531 -1121 -497
rect -1183 -537 -1121 -531
rect -1055 -497 -993 -491
rect -1055 -531 -1043 -497
rect -1005 -531 -993 -497
rect -1055 -537 -993 -531
rect -927 -497 -865 -491
rect -927 -531 -915 -497
rect -877 -531 -865 -497
rect -927 -537 -865 -531
rect -799 -497 -737 -491
rect -799 -531 -787 -497
rect -749 -531 -737 -497
rect -799 -537 -737 -531
rect -671 -497 -609 -491
rect -671 -531 -659 -497
rect -621 -531 -609 -497
rect -671 -537 -609 -531
rect -543 -497 -481 -491
rect -543 -531 -531 -497
rect -493 -531 -481 -497
rect -543 -537 -481 -531
rect -415 -497 -353 -491
rect -415 -531 -403 -497
rect -365 -531 -353 -497
rect -415 -537 -353 -531
rect -287 -497 -225 -491
rect -287 -531 -275 -497
rect -237 -531 -225 -497
rect -287 -537 -225 -531
rect -159 -497 -97 -491
rect -159 -531 -147 -497
rect -109 -531 -97 -497
rect -159 -537 -97 -531
rect -31 -497 31 -491
rect -31 -531 -19 -497
rect 19 -531 31 -497
rect -31 -537 31 -531
rect 97 -497 159 -491
rect 97 -531 109 -497
rect 147 -531 159 -497
rect 97 -537 159 -531
rect 225 -497 287 -491
rect 225 -531 237 -497
rect 275 -531 287 -497
rect 225 -537 287 -531
rect 353 -497 415 -491
rect 353 -531 365 -497
rect 403 -531 415 -497
rect 353 -537 415 -531
rect 481 -497 543 -491
rect 481 -531 493 -497
rect 531 -531 543 -497
rect 481 -537 543 -531
rect 609 -497 671 -491
rect 609 -531 621 -497
rect 659 -531 671 -497
rect 609 -537 671 -531
rect 737 -497 799 -491
rect 737 -531 749 -497
rect 787 -531 799 -497
rect 737 -537 799 -531
rect 865 -497 927 -491
rect 865 -531 877 -497
rect 915 -531 927 -497
rect 865 -537 927 -531
rect 993 -497 1055 -491
rect 993 -531 1005 -497
rect 1043 -531 1055 -497
rect 993 -537 1055 -531
rect 1121 -497 1183 -491
rect 1121 -531 1133 -497
rect 1171 -531 1183 -497
rect 1121 -537 1183 -531
rect 1249 -497 1311 -491
rect 1249 -531 1261 -497
rect 1299 -531 1311 -497
rect 1249 -537 1311 -531
<< properties >>
string FIXED_BBOX -1458 -616 1458 616
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 4.5 l 0.35 m 1 nf 21 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
