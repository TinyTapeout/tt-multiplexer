magic
tech sky130A
timestamp 1716279736
<< nwell >>
rect -1 -139 402 139
<< pwell >>
rect -1 139 402 266
rect -1 -266 402 -139
<< mvnmos >>
rect 140 173 190 215
rect 290 173 340 215
rect 140 -215 190 -173
rect 290 -215 340 -173
<< mvpmos >>
rect 61 64 111 106
rect 140 64 190 106
rect 219 64 269 106
rect 290 64 340 106
rect 61 -106 111 -64
rect 140 -106 190 -64
rect 219 -106 269 -64
rect 290 -106 340 -64
<< mvndiff >>
rect 111 211 140 215
rect 111 177 117 211
rect 134 177 140 211
rect 111 173 140 177
rect 190 211 290 215
rect 190 177 196 211
rect 284 177 290 211
rect 190 173 290 177
rect 340 211 369 215
rect 340 177 346 211
rect 363 177 369 211
rect 340 173 369 177
rect 111 -177 140 -173
rect 111 -211 117 -177
rect 134 -211 140 -177
rect 111 -215 140 -211
rect 190 -177 290 -173
rect 190 -211 196 -177
rect 284 -211 290 -177
rect 190 -215 290 -211
rect 340 -177 369 -173
rect 340 -211 346 -177
rect 363 -211 369 -177
rect 340 -215 369 -211
<< mvpdiff >>
rect 32 102 61 106
rect 32 68 38 102
rect 55 68 61 102
rect 32 64 61 68
rect 111 102 140 106
rect 111 68 117 102
rect 134 68 140 102
rect 111 64 140 68
rect 190 102 219 106
rect 190 68 196 102
rect 213 68 219 102
rect 190 64 219 68
rect 269 64 290 106
rect 340 102 369 106
rect 340 68 346 102
rect 363 68 369 102
rect 340 64 369 68
rect 32 -68 61 -64
rect 32 -102 38 -68
rect 55 -102 61 -68
rect 32 -106 61 -102
rect 111 -68 140 -64
rect 111 -102 117 -68
rect 134 -102 140 -68
rect 111 -106 140 -102
rect 190 -68 219 -64
rect 190 -102 196 -68
rect 213 -102 219 -68
rect 190 -106 219 -102
rect 269 -106 290 -64
rect 340 -68 369 -64
rect 340 -102 346 -68
rect 363 -102 369 -68
rect 340 -106 369 -102
<< mvndiffc >>
rect 117 177 134 211
rect 196 177 284 211
rect 346 177 363 211
rect 117 -211 134 -177
rect 196 -211 284 -177
rect 346 -211 363 -177
<< mvpdiffc >>
rect 38 68 55 102
rect 117 68 134 102
rect 196 68 213 102
rect 346 68 363 102
rect 38 -102 55 -68
rect 117 -102 134 -68
rect 196 -102 213 -68
rect 346 -102 363 -68
<< mvpsubdiff >>
rect 52 214 71 226
rect 52 197 53 214
rect 70 197 71 214
rect 52 185 71 197
rect 52 -197 71 -185
rect 52 -214 53 -197
rect 70 -214 71 -197
rect 52 -226 71 -214
<< mvnsubdiff >>
rect 32 -33 44 33
rect 252 -33 264 33
<< mvpsubdiffcont >>
rect 53 197 70 214
rect 53 -214 70 -197
<< mvnsubdiffcont >>
rect 44 -33 252 33
<< poly >>
rect 290 251 340 259
rect 290 234 295 251
rect 335 234 340 251
rect 140 215 190 228
rect 290 215 340 234
rect 140 165 190 173
rect 61 149 269 165
rect 290 160 340 173
rect 61 130 159 149
rect 261 130 269 149
rect 61 114 269 130
rect 61 106 111 114
rect 140 106 190 114
rect 219 106 269 114
rect 290 106 340 119
rect 61 51 111 64
rect 140 51 190 64
rect 219 51 269 64
rect 290 40 340 64
rect 290 23 295 40
rect 335 23 340 40
rect 290 15 340 23
rect 290 -23 340 -15
rect 290 -40 295 -23
rect 335 -40 340 -23
rect 61 -64 111 -51
rect 140 -64 190 -51
rect 219 -64 269 -51
rect 290 -64 340 -40
rect 61 -114 111 -106
rect 140 -114 190 -106
rect 219 -114 269 -106
rect 61 -130 269 -114
rect 290 -119 340 -106
rect 61 -149 159 -130
rect 261 -149 269 -130
rect 61 -165 269 -149
rect 140 -173 190 -165
rect 290 -173 340 -160
rect 140 -228 190 -215
rect 290 -234 340 -215
rect 290 -251 295 -234
rect 335 -251 340 -234
rect 290 -259 340 -251
<< polycont >>
rect 295 234 335 251
rect 159 130 261 149
rect 295 23 335 40
rect 295 -40 335 -23
rect 159 -149 261 -130
rect 295 -251 335 -234
<< locali >>
rect 287 234 293 251
rect 117 213 134 219
rect 188 208 196 211
rect 284 208 292 211
rect 188 180 194 208
rect 286 180 292 208
rect 188 177 196 180
rect 284 177 292 180
rect 338 177 346 211
rect 363 177 371 211
rect 38 104 55 110
rect 338 152 371 177
rect 151 149 371 152
rect 151 130 159 149
rect 261 148 371 149
rect 261 131 288 148
rect 342 131 371 148
rect 261 130 371 131
rect 151 127 371 130
rect 117 60 134 66
rect 196 104 213 110
rect 338 102 371 127
rect 338 68 346 102
rect 363 68 371 102
rect 38 33 55 51
rect 196 33 213 51
rect 36 10 44 33
rect 36 -10 41 10
rect 36 -33 44 -10
rect 252 -33 260 33
rect 335 23 343 40
rect 38 -51 55 -33
rect 196 -51 213 -33
rect 287 -40 295 -23
rect 38 -110 55 -104
rect 117 -66 134 -60
rect 196 -110 213 -104
rect 338 -102 346 -68
rect 363 -102 371 -68
rect 338 -127 371 -102
rect 151 -130 371 -127
rect 151 -149 159 -130
rect 261 -131 371 -130
rect 261 -148 288 -131
rect 342 -148 371 -131
rect 261 -149 371 -148
rect 151 -152 371 -149
rect 338 -177 371 -152
rect 188 -180 196 -177
rect 284 -180 292 -177
rect 188 -208 194 -180
rect 286 -208 292 -180
rect 188 -211 196 -208
rect 284 -211 292 -208
rect 338 -211 346 -177
rect 363 -211 371 -177
rect 117 -219 134 -213
rect 287 -251 293 -234
<< viali >>
rect 53 214 70 236
rect 293 234 295 251
rect 295 234 335 251
rect 335 234 346 251
rect 53 197 70 214
rect 53 183 70 197
rect 117 211 134 213
rect 117 177 134 211
rect 194 180 196 208
rect 196 180 284 208
rect 284 180 286 208
rect 38 102 55 104
rect 38 68 55 102
rect 38 51 55 68
rect 117 102 134 177
rect 288 131 342 148
rect 117 68 134 102
rect 117 66 134 68
rect 196 102 213 104
rect 196 68 213 102
rect 196 51 213 68
rect 41 -10 44 10
rect 44 -10 210 10
rect 282 23 295 40
rect 295 23 335 40
rect 38 -68 55 -51
rect 295 -40 335 -23
rect 335 -40 348 -23
rect 38 -102 55 -68
rect 38 -104 55 -102
rect 117 -68 134 -66
rect 117 -102 134 -68
rect 117 -177 134 -102
rect 196 -68 213 -51
rect 196 -102 213 -68
rect 196 -104 213 -102
rect 288 -148 342 -131
rect 53 -197 70 -183
rect 53 -214 70 -197
rect 53 -236 70 -214
rect 117 -211 134 -177
rect 194 -208 196 -180
rect 196 -208 284 -180
rect 284 -208 286 -180
rect 117 -213 134 -211
rect 293 -251 295 -234
rect 295 -251 335 -234
rect 335 -251 346 -234
<< metal1 >>
rect 50 236 240 257
rect 50 183 53 236
rect 70 234 240 236
rect 70 183 73 234
rect 50 177 73 183
rect 114 213 137 219
rect 35 104 58 110
rect 35 51 38 104
rect 55 51 58 104
rect 114 66 117 213
rect 134 66 137 213
rect 188 211 240 234
rect 287 251 352 254
rect 287 234 293 251
rect 346 234 352 251
rect 287 231 352 234
rect 188 208 292 211
rect 188 180 194 208
rect 286 180 292 208
rect 188 177 292 180
rect 282 148 379 151
rect 282 131 288 148
rect 342 131 379 148
rect 282 128 379 131
rect 114 60 137 66
rect 193 104 216 110
rect 35 44 58 51
rect 193 51 196 104
rect 213 51 216 104
rect 193 44 216 51
rect 35 10 216 44
rect 35 -10 41 10
rect 210 -10 216 10
rect 35 -44 216 -10
rect 35 -51 58 -44
rect 35 -104 38 -51
rect 55 -104 58 -51
rect 193 -51 216 -44
rect 35 -110 58 -104
rect 114 -66 137 -60
rect 50 -183 73 -177
rect 50 -236 53 -183
rect 70 -234 73 -183
rect 114 -213 117 -66
rect 134 -213 137 -66
rect 193 -104 196 -51
rect 213 -104 216 -51
rect 193 -110 216 -104
rect 252 40 341 43
rect 252 23 282 40
rect 335 23 341 40
rect 252 20 341 23
rect 252 -128 275 20
rect 355 -20 379 128
rect 289 -23 379 -20
rect 289 -40 295 -23
rect 348 -40 379 -23
rect 289 -43 379 -40
rect 252 -131 348 -128
rect 252 -148 288 -131
rect 342 -148 348 -131
rect 252 -151 348 -148
rect 114 -219 137 -213
rect 188 -180 292 -177
rect 188 -208 194 -180
rect 286 -208 292 -180
rect 188 -211 292 -208
rect 188 -234 240 -211
rect 70 -236 240 -234
rect 50 -257 240 -236
rect 287 -234 352 -231
rect 287 -251 293 -234
rect 346 -251 352 -234
rect 287 -254 352 -251
<< end >>
