magic
tech sky130A
magscale 1 2
timestamp 1718438769
<< nwell >>
rect 594 0 1827 470
<< pwell >>
rect 13 0 594 470
<< nmos >>
rect 160 263 510 293
rect 160 177 510 207
<< pmoshvt >>
rect 630 263 1680 293
rect 630 177 1680 207
<< ndiff >>
rect 160 338 510 346
rect 160 304 172 338
rect 498 304 510 338
rect 160 293 510 304
rect 160 252 510 263
rect 160 218 172 252
rect 498 218 510 252
rect 160 207 510 218
rect 160 166 510 177
rect 160 132 172 166
rect 498 132 510 166
rect 160 124 510 132
<< pdiff >>
rect 630 338 1680 346
rect 630 304 642 338
rect 1668 304 1680 338
rect 630 293 1680 304
rect 630 252 1680 263
rect 630 218 642 252
rect 1668 218 1680 252
rect 630 207 1680 218
rect 630 166 1680 177
rect 630 132 642 166
rect 1668 132 1680 166
rect 630 124 1680 132
<< ndiffc >>
rect 172 304 498 338
rect 172 218 498 252
rect 172 132 498 166
<< pdiffc >>
rect 642 304 1668 338
rect 642 218 1668 252
rect 642 132 1668 166
<< psubdiff >>
rect 72 400 136 434
rect 480 400 504 434
rect 72 370 106 400
rect 72 70 106 100
rect 72 36 136 70
rect 480 36 504 70
<< nsubdiff >>
rect 636 400 660 434
rect 1704 400 1768 434
rect 1734 370 1768 400
rect 1734 70 1768 100
rect 636 36 660 70
rect 1704 36 1768 70
<< psubdiffcont >>
rect 136 400 480 434
rect 72 100 106 370
rect 136 36 480 70
<< nsubdiffcont >>
rect 660 400 1704 434
rect 1734 100 1768 370
rect 660 36 1704 70
<< poly >>
rect 538 330 592 346
rect 538 293 548 330
rect 134 263 160 293
rect 510 263 548 293
rect 538 207 548 263
rect 134 177 160 207
rect 510 177 548 207
rect 538 140 548 177
rect 582 293 592 330
rect 582 263 630 293
rect 1680 263 1706 293
rect 582 207 592 263
rect 582 177 630 207
rect 1680 177 1706 207
rect 582 140 592 177
rect 538 124 592 140
<< polycont >>
rect 548 140 582 330
<< locali >>
rect 72 400 136 434
rect 480 400 510 434
rect 630 400 660 434
rect 1704 400 1768 434
rect 72 370 106 400
rect 1734 370 1768 400
rect 156 304 172 338
rect 498 304 514 338
rect 548 330 550 346
rect 156 218 172 252
rect 498 218 514 252
rect 156 132 172 166
rect 498 132 514 166
rect 548 124 550 140
rect 590 124 592 346
rect 626 304 642 338
rect 1668 304 1684 338
rect 626 218 642 252
rect 1668 218 1684 252
rect 626 132 642 166
rect 1668 132 1684 166
rect 72 70 106 100
rect 1734 70 1768 100
rect 72 36 136 70
rect 480 36 510 70
rect 630 36 660 70
rect 1704 36 1768 70
<< viali >>
rect 136 400 480 434
rect 660 400 1704 434
rect 72 100 106 370
rect 172 304 498 338
rect 550 330 590 346
rect 172 218 498 252
rect 172 132 498 166
rect 550 140 582 330
rect 582 140 590 330
rect 550 124 590 140
rect 642 304 1668 338
rect 642 218 1668 252
rect 642 132 1668 166
rect 1734 100 1768 370
rect 136 36 480 70
rect 660 36 1704 70
<< metal1 >>
rect 66 434 510 440
rect 66 400 136 434
rect 480 400 510 434
rect 66 394 510 400
rect 66 370 112 394
rect 66 100 72 370
rect 106 100 112 370
rect 160 338 510 394
rect 630 434 1774 440
rect 630 400 660 434
rect 1704 400 1774 434
rect 630 394 1774 400
rect 160 304 172 338
rect 498 304 510 338
rect 160 298 510 304
rect 544 352 596 358
rect 160 209 166 261
rect 504 209 510 261
rect 66 76 112 100
rect 160 166 510 172
rect 160 132 172 166
rect 498 132 510 166
rect 160 76 510 132
rect 630 338 1680 394
rect 630 304 642 338
rect 1668 304 1680 338
rect 630 298 1680 304
rect 1728 370 1774 394
rect 630 209 636 261
rect 1674 209 1680 261
rect 544 112 596 118
rect 630 166 1680 172
rect 630 132 642 166
rect 1668 132 1680 166
rect 66 70 510 76
rect 66 36 136 70
rect 480 36 510 70
rect 66 30 510 36
rect 630 76 1680 132
rect 1728 100 1734 370
rect 1768 100 1774 370
rect 1728 76 1774 100
rect 630 70 1774 76
rect 630 36 660 70
rect 1704 36 1774 70
rect 630 30 1774 36
<< via1 >>
rect 544 346 596 352
rect 166 252 504 261
rect 166 218 172 252
rect 172 218 498 252
rect 498 218 504 252
rect 166 209 504 218
rect 544 124 550 346
rect 550 124 590 346
rect 590 124 596 346
rect 636 252 1674 261
rect 636 218 642 252
rect 642 218 1668 252
rect 1668 218 1674 252
rect 636 209 1674 218
rect 544 118 596 124
<< metal2 >>
rect 458 392 682 444
rect 458 261 510 392
rect 160 209 166 261
rect 504 209 510 261
rect 544 352 596 358
rect 630 261 682 392
rect 630 209 636 261
rect 1674 209 1680 261
rect 544 0 596 118
<< properties >>
string FIXED_BBOX 0 0 1840 470
<< end >>
