/*
 * tt_defs.vh
 *
 * Shared defines
 *
 * Copyright (c) 2023 Sylvain Munaut <tnt@246tNt.com>
 * SPDX-License-Identifier: Apache-2.0
 */

`define TT_G_X  16
`define TT_G_Y  24

`define TT_N_IO 8
`define TT_N_O  8
`define TT_N_I  10
