VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_pg_1v8_4
  CLASS BLOCK ;
  FOREIGN tt_pg_1v8_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.200 BY 511.360 ;
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000 0.000 1.200 509.840 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.700 0.000 5.200 509.840 ;
    END
  END VPWR
  PIN GPWR
    DIRECTION OUTPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 5.700 0.000 9.200 509.840 ;
    END
  END GPWR
  PIN ctrl
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.200000 ;
    PORT
      LAYER met4 ;
        RECT 0.000 510.860 9.200 511.360 ;
    END
  END ctrl
  OBS
      LAYER nwell ;
        RECT 0.060 0.500 9.140 511.240 ;
      LAYER li1 ;
        RECT 0.190 0.630 9.010 511.060 ;
      LAYER met1 ;
        RECT 0.160 0.600 9.040 511.090 ;
      LAYER met2 ;
        RECT 0.160 1.010 9.040 511.240 ;
      LAYER met3 ;
        RECT 0.500 3.720 9.200 511.360 ;
      LAYER met4 ;
        RECT 2.675 510.340 3.025 510.460 ;
  END
END tt_pg_1v8_4
END LIBRARY

