magic
tech sky130A
magscale 1 2
timestamp 1718285775
<< metal1 >>
rect 54 21364 106 21370
rect 54 140 106 146
<< via1 >>
rect 166 22108 504 22250
rect 636 22108 1674 22250
rect 32 21462 190 21834
rect 1650 21462 1808 21834
rect 54 146 106 21364
<< metal2 >>
rect 542 22270 598 22280
rect 160 22108 166 22250
rect 504 22108 510 22250
rect 542 22140 598 22150
rect 630 22108 636 22250
rect 1674 22108 1680 22250
rect 32 21834 190 21840
rect 544 21758 596 21922
rect 1650 21834 1808 21840
rect 32 21456 190 21462
rect 222 21391 276 21706
rect 990 21538 1112 21656
rect 50 21370 106 21379
rect 138 21337 276 21391
rect 138 21237 192 21337
rect 994 21273 1112 21538
rect 1650 21456 1808 21462
rect 50 21221 54 21230
rect 54 140 106 146
<< via2 >>
rect 169 22113 391 22183
rect 542 22150 598 22270
rect 809 22113 1671 22173
rect 115 21465 185 21831
rect 50 21364 106 21370
rect 50 21230 54 21364
rect 54 21230 106 21364
rect 1655 21465 1725 21831
<< metal3 >>
rect 535 22274 605 22280
rect 535 22205 536 22274
rect 604 22205 605 22274
rect 110 22183 400 22188
rect 110 22113 169 22183
rect 391 22113 400 22183
rect 535 22150 542 22205
rect 598 22150 605 22205
rect 535 22140 605 22150
rect 800 22173 1680 22178
rect 110 22108 400 22113
rect 800 22113 809 22173
rect 1671 22113 1680 22173
rect 800 22108 1680 22113
rect 110 21994 190 22108
rect 800 22000 1040 22108
rect 110 21462 111 21994
rect 189 21840 190 21994
rect 340 21999 1040 22000
rect 340 21921 346 21999
rect 1034 21921 1040 21999
rect 340 21920 1040 21921
rect 189 21831 1730 21840
rect 189 21760 1655 21831
rect 189 21462 190 21760
rect 110 21456 190 21462
rect 1650 21465 1655 21760
rect 1725 21465 1730 21831
rect 1650 21456 1730 21465
rect 45 21374 1045 21375
rect 45 21370 341 21374
rect 45 21230 50 21370
rect 106 21230 341 21370
rect 45 21226 341 21230
rect 1039 21226 1045 21374
rect 45 21225 1045 21226
<< via3 >>
rect 536 22270 604 22274
rect 536 22205 542 22270
rect 542 22205 598 22270
rect 598 22205 604 22270
rect 111 21831 189 21994
rect 346 21921 1034 21999
rect 111 21465 115 21831
rect 115 21465 185 21831
rect 185 21465 189 21831
rect 111 21462 189 21465
rect 341 21226 1039 21374
<< metal4 >>
rect 0 22274 1840 22304
rect 0 22205 536 22274
rect 604 22205 1840 22274
rect 0 22204 1840 22205
rect 0 21994 240 22000
rect 0 21462 111 21994
rect 189 21462 240 21994
rect 0 0 240 21462
rect 340 21999 1040 22000
rect 340 21921 346 21999
rect 1034 21921 1040 21999
rect 340 21374 1040 21921
rect 340 21226 341 21374
rect 1039 21226 1040 21374
rect 340 0 1040 21226
rect 1140 0 1840 22000
use cap_gpwr  cap_gpwr_0
timestamp 1718097123
transform 1 0 0 0 1 3440
box 0 0 1840 4000
use cap_gpwr  cap_gpwr_1
timestamp 1718097123
transform 1 0 0 0 1 14864
box 0 0 1840 4000
use cap_vpwr  cap_vpwr_0
timestamp 1718097035
transform 1 0 0 0 1 9152
box 0 0 1840 4000
use ckt  ckt_0
timestamp 1718271279
transform 1 0 0 0 1 804
box 0 0 1840 1120
use ckt  ckt_1
timestamp 1718271279
transform 1 0 0 0 1 2024
box 0 0 1840 1120
use ckt  ckt_2
timestamp 1718271279
transform 1 0 0 0 1 7738
box 0 0 1840 1120
use ckt  ckt_3
timestamp 1718271279
transform 1 0 0 0 1 13448
box 0 0 1840 1120
use ckt  ckt_4
timestamp 1718271279
transform 1 0 0 0 1 19160
box 0 0 1840 1120
use discharge  discharge_0
timestamp 1718083762
transform 1 0 0 0 -1 21860
box 12 0 1828 424
use gate_inv  gate_inv_0
timestamp 1718283075
transform 1 0 0 0 -1 22280
box 13 0 1827 384
use pwr_pmos  pwr_pmos_0
timestamp 1718087245
transform -1 0 1810 0 1 110
box 0 0 1780 21290
<< labels >>
flabel metal4 s 0 0 240 22000 0 FreeSans 320 0 0 0 VGND
port 1 nsew ground input
flabel metal4 s 340 0 1040 22000 0 FreeSans 320 0 0 0 VPWR
port 2 nsew power input
flabel metal4 s 1140 0 1840 22000 0 FreeSans 320 0 0 0 GPWR
port 3 nsew power output
flabel metal4 s 0 22204 1840 22304 0 FreeSans 320 0 0 0 ctrl
port 4 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 1840 22304
<< end >>
