magic
tech sky130A
magscale 1 2
timestamp 1718543408
<< nwell >>
rect 1950 44030 2506 44246
rect 887 43210 2707 43360
<< metal1 >>
rect 332 45114 659 45148
rect 332 45038 366 45114
rect 593 45102 659 45114
rect 659 45052 2736 45098
rect 593 44954 659 44960
rect 2690 44952 2736 45052
rect 92 44822 1720 44868
rect 1790 44473 1796 44525
rect 2102 44473 2108 44525
rect 2348 44473 2354 44525
rect 2660 44473 2666 44525
rect 2617 43144 2669 43150
rect 2617 160 2669 166
<< via1 >>
rect 98 44960 270 45080
rect 426 44960 482 45080
rect 593 44960 659 45102
rect 20 44146 266 44658
rect 1406 44146 1652 44658
rect 1806 44630 1874 44826
rect 1796 44473 2102 44525
rect 2140 44324 2316 44674
rect 2582 44630 2650 44826
rect 2354 44473 2660 44525
rect 225 43828 813 43990
rect 959 43828 2547 43970
rect 225 43400 668 43562
rect 1104 43420 2547 43562
rect 2617 166 2669 43144
<< metal2 >>
rect 593 45102 659 45108
rect 92 45071 98 45080
rect 270 45071 276 45080
rect 92 44969 97 45071
rect 271 44969 276 45071
rect 92 44960 98 44969
rect 270 44960 276 44969
rect 420 45071 426 45080
rect 482 45071 488 45080
rect 593 44954 659 44960
rect 420 44926 488 44935
rect 1806 44826 1886 44832
rect 1874 44823 1886 44826
rect 1322 44708 1756 44760
rect 20 44658 266 44664
rect 1322 44562 1374 44708
rect 1406 44658 1652 44664
rect 906 44451 936 44460
rect 931 44251 936 44451
rect 906 44242 936 44251
rect 20 44140 266 44146
rect 1704 44525 1756 44708
rect 1881 44633 1886 44823
rect 2570 44826 2650 44832
rect 2570 44823 2582 44826
rect 1874 44630 1886 44633
rect 1806 44624 1886 44630
rect 2140 44674 2316 44680
rect 1704 44473 1796 44525
rect 2102 44473 2108 44525
rect 2570 44633 2575 44823
rect 2570 44630 2582 44633
rect 2570 44624 2650 44630
rect 2348 44473 2354 44525
rect 2660 44473 2666 44525
rect 2140 44318 2316 44324
rect 1406 44140 1652 44146
rect 2481 44082 2533 44473
rect 860 44030 2533 44082
rect 219 43828 225 43990
rect 813 43828 819 43990
rect 860 43876 912 44030
rect 953 43828 959 43970
rect 2547 43828 2553 43970
rect 219 43400 225 43562
rect 668 43400 674 43562
rect 1098 43420 1104 43562
rect 2547 43557 2669 43562
rect 2660 43487 2669 43557
rect 2547 43420 2669 43487
rect 715 43316 819 43358
rect 80 43212 819 43316
rect 80 42983 231 43212
rect 2617 43144 2669 43420
rect 80 327 177 42983
rect 2617 160 2669 166
<< via2 >>
rect 97 44969 98 45071
rect 98 44969 270 45071
rect 270 44969 271 45071
rect 420 44960 426 45071
rect 426 44960 482 45071
rect 482 44960 488 45071
rect 420 44935 488 44960
rect 598 44963 654 45099
rect 191 44149 261 44655
rect 771 44251 931 44451
rect 1411 44149 1481 44655
rect 1811 44633 1874 44823
rect 1874 44633 1881 44823
rect 2193 44327 2263 44671
rect 2575 44633 2582 44823
rect 2582 44633 2645 44823
rect 228 43833 727 43903
rect 1045 43833 2544 43903
rect 228 43487 665 43557
rect 1107 43487 2547 43557
rect 2547 43487 2660 43557
<< metal3 >>
rect 593 45146 659 45152
rect 26 45071 276 45080
rect 26 44969 97 45071
rect 271 44969 276 45071
rect 26 44960 276 44969
rect 414 45071 494 45080
rect 26 44847 106 44960
rect 26 44146 27 44847
rect 105 44146 106 44847
rect 414 44935 420 45071
rect 488 44935 494 45071
rect 593 44960 594 45146
rect 658 44960 659 45146
rect 593 44954 659 44960
rect 414 44664 494 44935
rect 1406 44823 2650 44832
rect 1406 44752 1811 44823
rect 1406 44664 1486 44752
rect 26 44140 106 44146
rect 186 44663 1486 44664
rect 186 44655 341 44663
rect 186 44149 191 44655
rect 261 44585 341 44655
rect 579 44655 1486 44663
rect 579 44585 1411 44655
rect 261 44584 1411 44585
rect 261 44149 266 44584
rect 766 44451 936 44460
rect 766 44251 771 44451
rect 931 44251 936 44451
rect 766 44242 936 44251
rect 186 43908 266 44149
rect 186 43907 736 43908
rect 186 43903 341 43907
rect 579 43903 736 43907
rect 186 43833 228 43903
rect 727 43833 736 43903
rect 186 43829 341 43833
rect 579 43829 736 43833
rect 186 43828 736 43829
rect 186 43562 266 43828
rect 186 43561 674 43562
rect 186 43557 341 43561
rect 579 43557 674 43561
rect 186 43487 228 43557
rect 665 43487 674 43557
rect 186 43483 341 43487
rect 579 43483 674 43487
rect 186 43482 674 43483
rect 836 43348 936 44242
rect 1406 44149 1411 44584
rect 1481 44149 1486 44655
rect 1806 44633 1811 44752
rect 1881 44752 2575 44823
rect 1881 44633 1886 44752
rect 1806 44624 1886 44633
rect 2188 44671 2268 44680
rect 1406 44140 1486 44149
rect 2188 44327 2193 44671
rect 2263 44327 2268 44671
rect 2570 44633 2575 44752
rect 2645 44633 2650 44823
rect 2570 44624 2650 44633
rect 2188 43908 2268 44327
rect 1036 43907 2553 43908
rect 1036 43829 1042 43907
rect 1669 43903 2553 43907
rect 2544 43833 2553 43903
rect 1669 43829 2553 43833
rect 1036 43828 2553 43829
rect 1098 43562 1178 43828
rect 1098 43561 2669 43562
rect 1098 43483 1104 43561
rect 1669 43557 2669 43561
rect 2660 43487 2669 43557
rect 1669 43483 2669 43487
rect 1098 43482 2669 43483
rect 836 43248 1724 43348
rect 1624 43128 1724 43248
<< via3 >>
rect 27 44146 105 44847
rect 594 45099 658 45146
rect 594 44963 598 45099
rect 598 44963 654 45099
rect 654 44963 658 45099
rect 594 44960 658 44963
rect 341 44585 579 44663
rect 341 43903 579 43907
rect 341 43833 579 43903
rect 341 43829 579 43833
rect 341 43557 579 43561
rect 341 43487 579 43557
rect 341 43483 579 43487
rect 1042 43903 1669 43907
rect 1042 43833 1045 43903
rect 1045 43833 1669 43903
rect 1042 43829 1669 43833
rect 1104 43557 1669 43561
rect 1104 43487 1107 43557
rect 1107 43487 1669 43557
rect 1104 43483 1669 43487
<< metal4 >>
rect 0 45146 2760 45152
rect 0 45052 594 45146
rect 593 44960 594 45052
rect 658 45052 2760 45146
rect 658 44960 659 45052
rect 593 44954 659 44960
rect 0 44847 240 44848
rect 0 44146 27 44847
rect 105 44146 240 44847
rect 0 0 240 44146
rect 340 44663 580 44848
rect 340 44585 341 44663
rect 579 44585 580 44663
rect 340 43907 580 44585
rect 340 43829 341 43907
rect 579 43829 580 43907
rect 340 43561 580 43829
rect 340 43483 341 43561
rect 579 43483 580 43561
rect 340 0 580 43483
rect 680 43907 1670 44848
rect 680 43829 1042 43907
rect 1669 43829 1670 43907
rect 680 43561 1670 43829
rect 680 43483 1104 43561
rect 1669 43483 1670 43561
rect 680 0 1670 43483
rect 1770 0 2760 44848
use cap_gapwr  cap_gapwr_0
timestamp 1718383489
transform 1 0 0 0 1 3440
box 0 0 2760 4000
use cap_gapwr  cap_gapwr_1
timestamp 1718383489
transform 1 0 0 0 1 14864
box 0 0 2760 4000
use cap_gapwr  cap_gapwr_2
timestamp 1718383489
transform 1 0 0 0 1 26288
box 0 0 2760 4000
use cap_gapwr  cap_gapwr_3
timestamp 1718383489
transform 1 0 0 0 1 37712
box 0 0 2760 4000
use cap_vapwr  cap_vapwr_0
timestamp 1718383489
transform 1 0 0 0 1 9152
box 0 0 2760 4000
use cap_vapwr  cap_vapwr_1
timestamp 1718383489
transform 1 0 0 0 1 32000
box 0 0 2760 4000
use ckt  ckt_0
timestamp 1718383489
transform 1 0 0 0 1 2024
box 0 0 2760 1120
use ckt  ckt_1
timestamp 1718383489
transform 1 0 0 0 1 7736
box 0 0 2760 1120
use ckt  ckt_2
timestamp 1718383489
transform 1 0 0 0 1 13448
box 0 0 2760 1120
use ckt  ckt_3
timestamp 1718383489
transform 1 0 0 0 1 19576
box 0 0 2760 1120
use ckt  ckt_4
timestamp 1718383489
transform 1 0 0 0 1 20796
box 0 0 2760 1120
use ckt  ckt_5
timestamp 1718383489
transform 1 0 0 0 1 22016
box 0 0 2760 1120
use ckt  ckt_6
timestamp 1718383489
transform 1 0 0 0 1 23236
box 0 0 2760 1120
use ckt  ckt_7
timestamp 1718383489
transform 1 0 0 0 1 24456
box 0 0 2760 1120
use ckt  ckt_8
timestamp 1718383489
transform 1 0 0 0 1 30584
box 0 0 2760 1120
use ckt  ckt_9
timestamp 1718383489
transform 1 0 0 0 1 36296
box 0 0 2760 1120
use ckt  ckt_10
timestamp 1718383489
transform 1 0 0 0 1 42008
box 0 0 2760 1120
use ctrl_inv  ctrl_inv_0
timestamp 1718543408
transform 0 1 -4796 -1 0 45770
box 668 4844 940 5328
use discharge  discharge_0
timestamp 1718532220
transform 1 0 0 0 -1 44684
box 0 0 1672 564
use gate_inv  gate_inv_0
timestamp 1718533623
transform 1 0 0 0 -1 44030
box 52 0 2707 672
use lv2hv  lv2hv_0
timestamp 1718383489
transform 0 1 2228 1 0 44248
box -2 -532 804 532
use pwr_pmos  pwr_pmos_0
timestamp 1718382556
transform 1 0 37 0 1 100
box 0 0 2686 43110
<< labels >>
flabel metal4 s 0 0 240 44848 0 FreeSans 320 0 0 0 VDPWR
port 1 nsew ground input
flabel metal4 s 340 0 580 44848 0 FreeSans 320 0 0 0 VGND
port 2 nsew ground input
flabel metal4 s 680 0 1670 44848 0 FreeSans 320 0 0 0 VAPWR
port 3 nsew power input
flabel metal4 s 1770 0 2760 44848 0 FreeSans 320 0 0 0 GAPWR
port 4 nsew power output
flabel metal4 s 0 45052 2760 45152 0 FreeSans 320 0 0 0 ctrl
port 5 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 2760 45152
<< end >>
