magic
tech sky130A
magscale 1 2
timestamp 1718289518
<< metal1 >>
rect 1734 100916 1786 100922
rect 1734 744 1786 750
<< via1 >>
rect 32 101070 190 101542
rect 1650 101070 1808 101542
rect 1734 750 1786 100916
<< metal2 >>
rect 542 102239 598 102248
rect 542 101716 598 101725
rect 32 101542 190 101548
rect 518 101466 624 101604
rect 1650 101542 1808 101548
rect 32 101064 190 101070
rect 518 100995 624 101414
rect 990 101146 1212 101364
rect 60 100889 624 100995
rect 60 100789 192 100889
rect 994 100825 1212 101146
rect 1650 101064 1808 101070
rect 1734 100917 1790 100926
rect 60 877 138 100789
rect 1786 100768 1790 100777
rect 1786 889 1790 898
rect 139 773 192 877
rect 139 720 275 773
rect 222 583 275 720
rect 222 254 274 583
rect 994 522 1212 841
rect 1734 740 1790 749
rect 990 304 1212 522
<< via2 >>
rect 119 102081 363 102151
rect 119 101701 363 101771
rect 542 101725 598 102239
rect 776 102081 1765 102151
rect 777 101701 1766 101771
rect 115 101073 185 101539
rect 1655 101073 1725 101539
rect 1734 100916 1790 100917
rect 1734 100777 1786 100916
rect 1786 100777 1790 100916
rect 1734 750 1786 889
rect 1786 750 1790 889
rect 1734 749 1790 750
<< metal3 >>
rect 535 102266 605 102272
rect 110 102151 372 102156
rect 110 102081 119 102151
rect 363 102081 372 102151
rect 110 102076 372 102081
rect 110 101962 190 102076
rect 110 101070 111 101962
rect 189 101776 190 101962
rect 535 102074 536 102266
rect 604 102074 605 102266
rect 189 101771 372 101776
rect 363 101701 372 101771
rect 535 101725 542 102074
rect 598 101725 605 102074
rect 535 101716 605 101725
rect 768 102151 1774 102156
rect 768 102081 776 102151
rect 1765 102081 1774 102151
rect 768 102076 1774 102081
rect 768 101824 848 102076
rect 768 101823 1040 101824
rect 189 101696 372 101701
rect 189 101460 190 101696
rect 768 101635 774 101823
rect 1034 101776 1040 101823
rect 1034 101771 1774 101776
rect 1766 101701 1774 101771
rect 1034 101696 1774 101701
rect 1034 101635 1040 101696
rect 768 101634 1040 101635
rect 1650 101539 1730 101548
rect 1650 101460 1655 101539
rect 189 101380 1655 101460
rect 189 101070 190 101380
rect 110 101064 190 101070
rect 1650 101073 1655 101380
rect 1725 101073 1730 101539
rect 1650 101064 1730 101073
rect 822 100921 1795 100922
rect 822 100773 828 100921
rect 1034 100917 1795 100921
rect 1034 100777 1734 100917
rect 1790 100777 1795 100917
rect 1034 100773 1795 100777
rect 822 100772 1795 100773
rect 822 893 1795 894
rect 822 745 828 893
rect 1034 889 1795 893
rect 1034 749 1734 889
rect 1790 749 1795 889
rect 1034 745 1795 749
rect 822 744 1795 745
<< via3 >>
rect 111 101771 189 101962
rect 536 102239 604 102266
rect 536 102074 542 102239
rect 542 102074 598 102239
rect 598 102074 604 102239
rect 111 101701 119 101771
rect 119 101701 189 101771
rect 111 101539 189 101701
rect 111 101073 115 101539
rect 115 101073 185 101539
rect 185 101073 189 101539
rect 774 101771 1034 101823
rect 774 101701 777 101771
rect 777 101701 1034 101771
rect 774 101635 1034 101701
rect 111 101070 189 101073
rect 828 100773 1034 100921
rect 828 745 1034 893
<< metal4 >>
rect 0 102266 1840 102272
rect 0 102172 536 102266
rect 535 102074 536 102172
rect 604 102172 1840 102266
rect 604 102074 605 102172
rect 535 102068 605 102074
rect 0 101962 240 101968
rect 0 101070 111 101962
rect 189 101070 240 101962
rect 0 0 240 101070
rect 340 101823 1040 101968
rect 340 101635 774 101823
rect 1034 101635 1040 101823
rect 340 100921 1040 101635
rect 340 100773 828 100921
rect 1034 100773 1040 100921
rect 340 893 1040 100773
rect 340 745 828 893
rect 1034 745 1040 893
rect 340 0 1040 745
rect 1140 0 1840 101968
use cap_gpwr  cap_gpwr_0
timestamp 1718097123
transform 1 0 0 0 1 3440
box 0 0 1840 4000
use cap_gpwr  cap_gpwr_1
timestamp 1718097123
transform 1 0 0 0 1 14864
box 0 0 1840 4000
use cap_gpwr  cap_gpwr_3
timestamp 1718097123
transform 1 0 0 0 1 26288
box 0 0 1840 4000
use cap_gpwr  cap_gpwr_4
timestamp 1718097123
transform 1 0 0 0 1 37712
box 0 0 1840 4000
use cap_gpwr  cap_gpwr_5
timestamp 1718097123
transform 1 0 0 0 1 49136
box 0 0 1840 4000
use cap_gpwr  cap_gpwr_6
timestamp 1718097123
transform 1 0 0 0 1 60560
box 0 0 1840 4000
use cap_gpwr  cap_gpwr_7
timestamp 1718097123
transform 1 0 0 0 1 71984
box 0 0 1840 4000
use cap_gpwr  cap_gpwr_8
timestamp 1718097123
transform 1 0 0 0 1 83408
box 0 0 1840 4000
use cap_gpwr  cap_gpwr_9
timestamp 1718097123
transform 1 0 0 0 1 94832
box 0 0 1840 4000
use cap_vpwr  cap_vpwr_0
timestamp 1718097035
transform 1 0 0 0 1 9152
box 0 0 1840 4000
use cap_vpwr  cap_vpwr_1
timestamp 1718097035
transform 1 0 0 0 1 89120
box 0 0 1840 4000
use cap_vpwr  cap_vpwr_2
timestamp 1718097035
transform 1 0 0 0 1 20576
box 0 0 1840 4000
use cap_vpwr  cap_vpwr_3
timestamp 1718097035
transform 1 0 0 0 1 43424
box 0 0 1840 4000
use cap_vpwr  cap_vpwr_4
timestamp 1718097035
transform 1 0 0 0 1 54848
box 0 0 1840 4000
use cap_vpwr  cap_vpwr_5
timestamp 1718097035
transform 1 0 0 0 1 77696
box 0 0 1840 4000
use ckt  ckt_0
timestamp 1718271279
transform 1 0 0 0 1 2024
box 0 0 1840 1120
use ckt  ckt_1
timestamp 1718271279
transform 1 0 0 0 1 7736
box 0 0 1840 1120
use ckt  ckt_2
timestamp 1718271279
transform 1 0 0 0 1 13448
box 0 0 1840 1120
use ckt  ckt_3
timestamp 1718271279
transform 1 0 0 0 1 19160
box 0 0 1840 1120
use ckt  ckt_4
timestamp 1718271279
transform 1 0 0 0 1 24872
box 0 0 1840 1120
use ckt  ckt_5
timestamp 1718271279
transform 1 0 0 0 1 30950
box 0 0 1840 1120
use ckt  ckt_6
timestamp 1718271279
transform 1 0 0 0 1 32170
box 0 0 1840 1120
use ckt  ckt_7
timestamp 1718271279
transform 1 0 0 0 1 33390
box 0 0 1840 1120
use ckt  ckt_8
timestamp 1718271279
transform 1 0 0 0 1 34610
box 0 0 1840 1120
use ckt  ckt_9
timestamp 1718271279
transform 1 0 0 0 1 35830
box 0 0 1840 1120
use ckt  ckt_10
timestamp 1718271279
transform 1 0 0 0 1 42008
box 0 0 1840 1120
use ckt  ckt_11
timestamp 1718271279
transform 1 0 0 0 1 47720
box 0 0 1840 1120
use ckt  ckt_12
timestamp 1718271279
transform 1 0 0 0 1 53432
box 0 0 1840 1120
use ckt  ckt_13
timestamp 1718271279
transform 1 0 0 0 1 59144
box 0 0 1840 1120
use ckt  ckt_14
timestamp 1718271279
transform 1 0 0 0 1 65222
box 0 0 1840 1120
use ckt  ckt_15
timestamp 1718271279
transform 1 0 0 0 1 66442
box 0 0 1840 1120
use ckt  ckt_16
timestamp 1718271279
transform 1 0 0 0 1 67662
box 0 0 1840 1120
use ckt  ckt_17
timestamp 1718271279
transform 1 0 0 0 1 68882
box 0 0 1840 1120
use ckt  ckt_18
timestamp 1718271279
transform 1 0 0 0 1 70102
box 0 0 1840 1120
use ckt  ckt_19
timestamp 1718271279
transform 1 0 0 0 1 76280
box 0 0 1840 1120
use ckt  ckt_20
timestamp 1718271279
transform 1 0 0 0 1 81992
box 0 0 1840 1120
use ckt  ckt_21
timestamp 1718271279
transform 1 0 0 0 1 87704
box 0 0 1840 1120
use ckt  ckt_22
timestamp 1718271279
transform 1 0 0 0 1 93416
box 0 0 1840 1120
use ckt  ckt_23
timestamp 1718271279
transform 1 0 0 0 1 99128
box 0 0 1840 1120
use discharge  discharge_0
timestamp 1718199492
transform 1 0 0 0 1 100
box 12 0 1828 524
use discharge  discharge_1
timestamp 1718199492
transform 1 0 0 0 -1 101568
box 12 0 1828 524
use gate_inv  gate_inv_0
timestamp 1718283606
transform 1 0 0 0 -1 102248
box 13 0 1827 644
use pwr_pmos  pwr_pmos_0
timestamp 1718224900
transform -1 0 1810 0 1 714
box 0 0 1780 100238
<< labels >>
flabel metal4 s 0 0 240 101968 0 FreeSans 320 0 0 0 VGND
port 1 nsew ground input
flabel metal4 s 340 0 1040 101968 0 FreeSans 320 0 0 0 VPWR
port 2 nsew power input
flabel metal4 s 1140 0 1840 101968 0 FreeSans 320 0 0 0 GPWR
port 3 nsew power output
flabel metal4 s 0 102172 1840 102272 0 FreeSans 320 0 0 0 ctrl
port 4 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 1840 102272
<< end >>
