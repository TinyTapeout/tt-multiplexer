VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO vccd1_connection
  CLASS BLOCK ;
  FOREIGN vccd1_connection ;
  ORIGIN 0.000 0.000 ;
  SIZE 45.400 BY 74.600 ;
  OBS
      LAYER met3 ;
        RECT 0.105 0.100 45.340 74.300 ;
  END
END vccd1_connection
END LIBRARY

