magic
tech sky130A
magscale 1 2
timestamp 1718224900
<< nwell >>
rect 0 0 1780 100238
<< pmos >>
rect 130 100027 1580 100057
rect 130 99941 1580 99971
rect 130 99855 1580 99885
rect 130 99769 1580 99799
rect 130 99683 1580 99713
rect 130 99597 1580 99627
rect 130 99511 1580 99541
rect 130 99425 1580 99455
rect 130 99339 1580 99369
rect 130 99253 1580 99283
rect 130 99167 1580 99197
rect 130 99081 1580 99111
rect 130 98995 1580 99025
rect 130 98909 1580 98939
rect 130 98823 1580 98853
rect 130 98737 1580 98767
rect 130 98651 1580 98681
rect 130 98565 1580 98595
rect 130 98479 1580 98509
rect 130 98393 1580 98423
rect 130 98307 1580 98337
rect 130 98221 1580 98251
rect 130 98135 1580 98165
rect 130 98049 1580 98079
rect 130 97963 1580 97993
rect 130 97877 1580 97907
rect 130 97791 1580 97821
rect 130 97705 1580 97735
rect 130 97619 1580 97649
rect 130 97533 1580 97563
rect 130 97447 1580 97477
rect 130 97361 1580 97391
rect 130 97275 1580 97305
rect 130 97189 1580 97219
rect 130 97103 1580 97133
rect 130 97017 1580 97047
rect 130 96931 1580 96961
rect 130 96845 1580 96875
rect 130 96759 1580 96789
rect 130 96673 1580 96703
rect 130 96587 1580 96617
rect 130 96501 1580 96531
rect 130 96415 1580 96445
rect 130 96329 1580 96359
rect 130 96243 1580 96273
rect 130 96157 1580 96187
rect 130 96071 1580 96101
rect 130 95985 1580 96015
rect 130 95899 1580 95929
rect 130 95813 1580 95843
rect 130 95727 1580 95757
rect 130 95641 1580 95671
rect 130 95555 1580 95585
rect 130 95469 1580 95499
rect 130 95383 1580 95413
rect 130 95297 1580 95327
rect 130 95211 1580 95241
rect 130 95125 1580 95155
rect 130 95039 1580 95069
rect 130 94953 1580 94983
rect 130 94867 1580 94897
rect 130 94781 1580 94811
rect 130 94695 1580 94725
rect 130 94609 1580 94639
rect 130 94523 1580 94553
rect 130 94437 1580 94467
rect 130 94351 1580 94381
rect 130 94265 1580 94295
rect 130 94179 1580 94209
rect 130 94093 1580 94123
rect 130 94007 1580 94037
rect 130 93921 1580 93951
rect 130 93835 1580 93865
rect 130 93749 1580 93779
rect 130 93663 1580 93693
rect 130 93577 1580 93607
rect 130 93491 1580 93521
rect 130 93405 1580 93435
rect 130 93319 1580 93349
rect 130 93233 1580 93263
rect 130 93147 1580 93177
rect 130 93061 1580 93091
rect 130 92975 1580 93005
rect 130 92889 1580 92919
rect 130 92803 1580 92833
rect 130 92717 1580 92747
rect 130 92631 1580 92661
rect 130 92545 1580 92575
rect 130 92459 1580 92489
rect 130 92373 1580 92403
rect 130 92287 1580 92317
rect 130 92201 1580 92231
rect 130 92115 1580 92145
rect 130 92029 1580 92059
rect 130 91943 1580 91973
rect 130 91857 1580 91887
rect 130 91771 1580 91801
rect 130 91685 1580 91715
rect 130 91599 1580 91629
rect 130 91513 1580 91543
rect 130 91427 1580 91457
rect 130 91341 1580 91371
rect 130 91255 1580 91285
rect 130 91169 1580 91199
rect 130 91083 1580 91113
rect 130 90997 1580 91027
rect 130 90911 1580 90941
rect 130 90825 1580 90855
rect 130 90739 1580 90769
rect 130 90653 1580 90683
rect 130 90567 1580 90597
rect 130 90481 1580 90511
rect 130 90395 1580 90425
rect 130 90309 1580 90339
rect 130 90223 1580 90253
rect 130 90137 1580 90167
rect 130 90051 1580 90081
rect 130 89965 1580 89995
rect 130 89879 1580 89909
rect 130 89793 1580 89823
rect 130 89707 1580 89737
rect 130 89621 1580 89651
rect 130 89535 1580 89565
rect 130 89449 1580 89479
rect 130 89363 1580 89393
rect 130 89277 1580 89307
rect 130 89191 1580 89221
rect 130 89105 1580 89135
rect 130 89019 1580 89049
rect 130 88933 1580 88963
rect 130 88847 1580 88877
rect 130 88761 1580 88791
rect 130 88675 1580 88705
rect 130 88589 1580 88619
rect 130 88503 1580 88533
rect 130 88417 1580 88447
rect 130 88331 1580 88361
rect 130 88245 1580 88275
rect 130 88159 1580 88189
rect 130 88073 1580 88103
rect 130 87987 1580 88017
rect 130 87901 1580 87931
rect 130 87815 1580 87845
rect 130 87729 1580 87759
rect 130 87643 1580 87673
rect 130 87557 1580 87587
rect 130 87471 1580 87501
rect 130 87385 1580 87415
rect 130 87299 1580 87329
rect 130 87213 1580 87243
rect 130 87127 1580 87157
rect 130 87041 1580 87071
rect 130 86955 1580 86985
rect 130 86869 1580 86899
rect 130 86783 1580 86813
rect 130 86697 1580 86727
rect 130 86611 1580 86641
rect 130 86525 1580 86555
rect 130 86439 1580 86469
rect 130 86353 1580 86383
rect 130 86267 1580 86297
rect 130 86181 1580 86211
rect 130 86095 1580 86125
rect 130 86009 1580 86039
rect 130 85923 1580 85953
rect 130 85837 1580 85867
rect 130 85751 1580 85781
rect 130 85665 1580 85695
rect 130 85579 1580 85609
rect 130 85493 1580 85523
rect 130 85407 1580 85437
rect 130 85321 1580 85351
rect 130 85235 1580 85265
rect 130 85149 1580 85179
rect 130 85063 1580 85093
rect 130 84977 1580 85007
rect 130 84891 1580 84921
rect 130 84805 1580 84835
rect 130 84719 1580 84749
rect 130 84633 1580 84663
rect 130 84547 1580 84577
rect 130 84461 1580 84491
rect 130 84375 1580 84405
rect 130 84289 1580 84319
rect 130 84203 1580 84233
rect 130 84117 1580 84147
rect 130 84031 1580 84061
rect 130 83945 1580 83975
rect 130 83859 1580 83889
rect 130 83773 1580 83803
rect 130 83687 1580 83717
rect 130 83601 1580 83631
rect 130 83515 1580 83545
rect 130 83429 1580 83459
rect 130 83343 1580 83373
rect 130 83257 1580 83287
rect 130 83171 1580 83201
rect 130 83085 1580 83115
rect 130 82999 1580 83029
rect 130 82913 1580 82943
rect 130 82827 1580 82857
rect 130 82741 1580 82771
rect 130 82655 1580 82685
rect 130 82569 1580 82599
rect 130 82483 1580 82513
rect 130 82397 1580 82427
rect 130 82311 1580 82341
rect 130 82225 1580 82255
rect 130 82139 1580 82169
rect 130 82053 1580 82083
rect 130 81967 1580 81997
rect 130 81881 1580 81911
rect 130 81795 1580 81825
rect 130 81709 1580 81739
rect 130 81623 1580 81653
rect 130 81537 1580 81567
rect 130 81451 1580 81481
rect 130 81365 1580 81395
rect 130 81279 1580 81309
rect 130 81193 1580 81223
rect 130 81107 1580 81137
rect 130 81021 1580 81051
rect 130 80935 1580 80965
rect 130 80849 1580 80879
rect 130 80763 1580 80793
rect 130 80677 1580 80707
rect 130 80591 1580 80621
rect 130 80505 1580 80535
rect 130 80419 1580 80449
rect 130 80333 1580 80363
rect 130 80247 1580 80277
rect 130 80161 1580 80191
rect 130 80075 1580 80105
rect 130 79989 1580 80019
rect 130 79903 1580 79933
rect 130 79817 1580 79847
rect 130 79731 1580 79761
rect 130 79645 1580 79675
rect 130 79559 1580 79589
rect 130 79473 1580 79503
rect 130 79387 1580 79417
rect 130 79301 1580 79331
rect 130 79215 1580 79245
rect 130 79129 1580 79159
rect 130 79043 1580 79073
rect 130 78957 1580 78987
rect 130 78871 1580 78901
rect 130 78785 1580 78815
rect 130 78699 1580 78729
rect 130 78613 1580 78643
rect 130 78527 1580 78557
rect 130 78441 1580 78471
rect 130 78355 1580 78385
rect 130 78269 1580 78299
rect 130 78183 1580 78213
rect 130 78097 1580 78127
rect 130 78011 1580 78041
rect 130 77925 1580 77955
rect 130 77839 1580 77869
rect 130 77753 1580 77783
rect 130 77667 1580 77697
rect 130 77581 1580 77611
rect 130 77495 1580 77525
rect 130 77409 1580 77439
rect 130 77323 1580 77353
rect 130 77237 1580 77267
rect 130 77151 1580 77181
rect 130 77065 1580 77095
rect 130 76979 1580 77009
rect 130 76893 1580 76923
rect 130 76807 1580 76837
rect 130 76721 1580 76751
rect 130 76635 1580 76665
rect 130 76549 1580 76579
rect 130 76463 1580 76493
rect 130 76377 1580 76407
rect 130 76291 1580 76321
rect 130 76205 1580 76235
rect 130 76119 1580 76149
rect 130 76033 1580 76063
rect 130 75947 1580 75977
rect 130 75861 1580 75891
rect 130 75775 1580 75805
rect 130 75689 1580 75719
rect 130 75603 1580 75633
rect 130 75517 1580 75547
rect 130 75431 1580 75461
rect 130 75345 1580 75375
rect 130 75259 1580 75289
rect 130 75173 1580 75203
rect 130 75087 1580 75117
rect 130 75001 1580 75031
rect 130 74915 1580 74945
rect 130 74829 1580 74859
rect 130 74743 1580 74773
rect 130 74657 1580 74687
rect 130 74571 1580 74601
rect 130 74485 1580 74515
rect 130 74399 1580 74429
rect 130 74313 1580 74343
rect 130 74227 1580 74257
rect 130 74141 1580 74171
rect 130 74055 1580 74085
rect 130 73969 1580 73999
rect 130 73883 1580 73913
rect 130 73797 1580 73827
rect 130 73711 1580 73741
rect 130 73625 1580 73655
rect 130 73539 1580 73569
rect 130 73453 1580 73483
rect 130 73367 1580 73397
rect 130 73281 1580 73311
rect 130 73195 1580 73225
rect 130 73109 1580 73139
rect 130 73023 1580 73053
rect 130 72937 1580 72967
rect 130 72851 1580 72881
rect 130 72765 1580 72795
rect 130 72679 1580 72709
rect 130 72593 1580 72623
rect 130 72507 1580 72537
rect 130 72421 1580 72451
rect 130 72335 1580 72365
rect 130 72249 1580 72279
rect 130 72163 1580 72193
rect 130 72077 1580 72107
rect 130 71991 1580 72021
rect 130 71905 1580 71935
rect 130 71819 1580 71849
rect 130 71733 1580 71763
rect 130 71647 1580 71677
rect 130 71561 1580 71591
rect 130 71475 1580 71505
rect 130 71389 1580 71419
rect 130 71303 1580 71333
rect 130 71217 1580 71247
rect 130 71131 1580 71161
rect 130 71045 1580 71075
rect 130 70959 1580 70989
rect 130 70873 1580 70903
rect 130 70787 1580 70817
rect 130 70701 1580 70731
rect 130 70615 1580 70645
rect 130 70529 1580 70559
rect 130 70443 1580 70473
rect 130 70357 1580 70387
rect 130 70271 1580 70301
rect 130 70185 1580 70215
rect 130 70099 1580 70129
rect 130 70013 1580 70043
rect 130 69927 1580 69957
rect 130 69841 1580 69871
rect 130 69755 1580 69785
rect 130 69669 1580 69699
rect 130 69583 1580 69613
rect 130 69497 1580 69527
rect 130 69411 1580 69441
rect 130 69325 1580 69355
rect 130 69239 1580 69269
rect 130 69153 1580 69183
rect 130 69067 1580 69097
rect 130 68981 1580 69011
rect 130 68895 1580 68925
rect 130 68809 1580 68839
rect 130 68723 1580 68753
rect 130 68637 1580 68667
rect 130 68551 1580 68581
rect 130 68465 1580 68495
rect 130 68379 1580 68409
rect 130 68293 1580 68323
rect 130 68207 1580 68237
rect 130 68121 1580 68151
rect 130 68035 1580 68065
rect 130 67949 1580 67979
rect 130 67863 1580 67893
rect 130 67777 1580 67807
rect 130 67691 1580 67721
rect 130 67605 1580 67635
rect 130 67519 1580 67549
rect 130 67433 1580 67463
rect 130 67347 1580 67377
rect 130 67261 1580 67291
rect 130 67175 1580 67205
rect 130 67089 1580 67119
rect 130 67003 1580 67033
rect 130 66917 1580 66947
rect 130 66831 1580 66861
rect 130 66745 1580 66775
rect 130 66659 1580 66689
rect 130 66573 1580 66603
rect 130 66487 1580 66517
rect 130 66401 1580 66431
rect 130 66315 1580 66345
rect 130 66229 1580 66259
rect 130 66143 1580 66173
rect 130 66057 1580 66087
rect 130 65971 1580 66001
rect 130 65885 1580 65915
rect 130 65799 1580 65829
rect 130 65713 1580 65743
rect 130 65627 1580 65657
rect 130 65541 1580 65571
rect 130 65455 1580 65485
rect 130 65369 1580 65399
rect 130 65283 1580 65313
rect 130 65197 1580 65227
rect 130 65111 1580 65141
rect 130 65025 1580 65055
rect 130 64939 1580 64969
rect 130 64853 1580 64883
rect 130 64767 1580 64797
rect 130 64681 1580 64711
rect 130 64595 1580 64625
rect 130 64509 1580 64539
rect 130 64423 1580 64453
rect 130 64337 1580 64367
rect 130 64251 1580 64281
rect 130 64165 1580 64195
rect 130 64079 1580 64109
rect 130 63993 1580 64023
rect 130 63907 1580 63937
rect 130 63821 1580 63851
rect 130 63735 1580 63765
rect 130 63649 1580 63679
rect 130 63563 1580 63593
rect 130 63477 1580 63507
rect 130 63391 1580 63421
rect 130 63305 1580 63335
rect 130 63219 1580 63249
rect 130 63133 1580 63163
rect 130 63047 1580 63077
rect 130 62961 1580 62991
rect 130 62875 1580 62905
rect 130 62789 1580 62819
rect 130 62703 1580 62733
rect 130 62617 1580 62647
rect 130 62531 1580 62561
rect 130 62445 1580 62475
rect 130 62359 1580 62389
rect 130 62273 1580 62303
rect 130 62187 1580 62217
rect 130 62101 1580 62131
rect 130 62015 1580 62045
rect 130 61929 1580 61959
rect 130 61843 1580 61873
rect 130 61757 1580 61787
rect 130 61671 1580 61701
rect 130 61585 1580 61615
rect 130 61499 1580 61529
rect 130 61413 1580 61443
rect 130 61327 1580 61357
rect 130 61241 1580 61271
rect 130 61155 1580 61185
rect 130 61069 1580 61099
rect 130 60983 1580 61013
rect 130 60897 1580 60927
rect 130 60811 1580 60841
rect 130 60725 1580 60755
rect 130 60639 1580 60669
rect 130 60553 1580 60583
rect 130 60467 1580 60497
rect 130 60381 1580 60411
rect 130 60295 1580 60325
rect 130 60209 1580 60239
rect 130 60123 1580 60153
rect 130 60037 1580 60067
rect 130 59951 1580 59981
rect 130 59865 1580 59895
rect 130 59779 1580 59809
rect 130 59693 1580 59723
rect 130 59607 1580 59637
rect 130 59521 1580 59551
rect 130 59435 1580 59465
rect 130 59349 1580 59379
rect 130 59263 1580 59293
rect 130 59177 1580 59207
rect 130 59091 1580 59121
rect 130 59005 1580 59035
rect 130 58919 1580 58949
rect 130 58833 1580 58863
rect 130 58747 1580 58777
rect 130 58661 1580 58691
rect 130 58575 1580 58605
rect 130 58489 1580 58519
rect 130 58403 1580 58433
rect 130 58317 1580 58347
rect 130 58231 1580 58261
rect 130 58145 1580 58175
rect 130 58059 1580 58089
rect 130 57973 1580 58003
rect 130 57887 1580 57917
rect 130 57801 1580 57831
rect 130 57715 1580 57745
rect 130 57629 1580 57659
rect 130 57543 1580 57573
rect 130 57457 1580 57487
rect 130 57371 1580 57401
rect 130 57285 1580 57315
rect 130 57199 1580 57229
rect 130 57113 1580 57143
rect 130 57027 1580 57057
rect 130 56941 1580 56971
rect 130 56855 1580 56885
rect 130 56769 1580 56799
rect 130 56683 1580 56713
rect 130 56597 1580 56627
rect 130 56511 1580 56541
rect 130 56425 1580 56455
rect 130 56339 1580 56369
rect 130 56253 1580 56283
rect 130 56167 1580 56197
rect 130 56081 1580 56111
rect 130 55995 1580 56025
rect 130 55909 1580 55939
rect 130 55823 1580 55853
rect 130 55737 1580 55767
rect 130 55651 1580 55681
rect 130 55565 1580 55595
rect 130 55479 1580 55509
rect 130 55393 1580 55423
rect 130 55307 1580 55337
rect 130 55221 1580 55251
rect 130 55135 1580 55165
rect 130 55049 1580 55079
rect 130 54963 1580 54993
rect 130 54877 1580 54907
rect 130 54791 1580 54821
rect 130 54705 1580 54735
rect 130 54619 1580 54649
rect 130 54533 1580 54563
rect 130 54447 1580 54477
rect 130 54361 1580 54391
rect 130 54275 1580 54305
rect 130 54189 1580 54219
rect 130 54103 1580 54133
rect 130 54017 1580 54047
rect 130 53931 1580 53961
rect 130 53845 1580 53875
rect 130 53759 1580 53789
rect 130 53673 1580 53703
rect 130 53587 1580 53617
rect 130 53501 1580 53531
rect 130 53415 1580 53445
rect 130 53329 1580 53359
rect 130 53243 1580 53273
rect 130 53157 1580 53187
rect 130 53071 1580 53101
rect 130 52985 1580 53015
rect 130 52899 1580 52929
rect 130 52813 1580 52843
rect 130 52727 1580 52757
rect 130 52641 1580 52671
rect 130 52555 1580 52585
rect 130 52469 1580 52499
rect 130 52383 1580 52413
rect 130 52297 1580 52327
rect 130 52211 1580 52241
rect 130 52125 1580 52155
rect 130 52039 1580 52069
rect 130 51953 1580 51983
rect 130 51867 1580 51897
rect 130 51781 1580 51811
rect 130 51695 1580 51725
rect 130 51609 1580 51639
rect 130 51523 1580 51553
rect 130 51437 1580 51467
rect 130 51351 1580 51381
rect 130 51265 1580 51295
rect 130 51179 1580 51209
rect 130 51093 1580 51123
rect 130 51007 1580 51037
rect 130 50921 1580 50951
rect 130 50835 1580 50865
rect 130 50749 1580 50779
rect 130 50663 1580 50693
rect 130 50577 1580 50607
rect 130 50491 1580 50521
rect 130 50405 1580 50435
rect 130 50319 1580 50349
rect 130 50233 1580 50263
rect 130 50147 1580 50177
rect 130 50061 1580 50091
rect 130 49975 1580 50005
rect 130 49889 1580 49919
rect 130 49803 1580 49833
rect 130 49717 1580 49747
rect 130 49631 1580 49661
rect 130 49545 1580 49575
rect 130 49459 1580 49489
rect 130 49373 1580 49403
rect 130 49287 1580 49317
rect 130 49201 1580 49231
rect 130 49115 1580 49145
rect 130 49029 1580 49059
rect 130 48943 1580 48973
rect 130 48857 1580 48887
rect 130 48771 1580 48801
rect 130 48685 1580 48715
rect 130 48599 1580 48629
rect 130 48513 1580 48543
rect 130 48427 1580 48457
rect 130 48341 1580 48371
rect 130 48255 1580 48285
rect 130 48169 1580 48199
rect 130 48083 1580 48113
rect 130 47997 1580 48027
rect 130 47911 1580 47941
rect 130 47825 1580 47855
rect 130 47739 1580 47769
rect 130 47653 1580 47683
rect 130 47567 1580 47597
rect 130 47481 1580 47511
rect 130 47395 1580 47425
rect 130 47309 1580 47339
rect 130 47223 1580 47253
rect 130 47137 1580 47167
rect 130 47051 1580 47081
rect 130 46965 1580 46995
rect 130 46879 1580 46909
rect 130 46793 1580 46823
rect 130 46707 1580 46737
rect 130 46621 1580 46651
rect 130 46535 1580 46565
rect 130 46449 1580 46479
rect 130 46363 1580 46393
rect 130 46277 1580 46307
rect 130 46191 1580 46221
rect 130 46105 1580 46135
rect 130 46019 1580 46049
rect 130 45933 1580 45963
rect 130 45847 1580 45877
rect 130 45761 1580 45791
rect 130 45675 1580 45705
rect 130 45589 1580 45619
rect 130 45503 1580 45533
rect 130 45417 1580 45447
rect 130 45331 1580 45361
rect 130 45245 1580 45275
rect 130 45159 1580 45189
rect 130 45073 1580 45103
rect 130 44987 1580 45017
rect 130 44901 1580 44931
rect 130 44815 1580 44845
rect 130 44729 1580 44759
rect 130 44643 1580 44673
rect 130 44557 1580 44587
rect 130 44471 1580 44501
rect 130 44385 1580 44415
rect 130 44299 1580 44329
rect 130 44213 1580 44243
rect 130 44127 1580 44157
rect 130 44041 1580 44071
rect 130 43955 1580 43985
rect 130 43869 1580 43899
rect 130 43783 1580 43813
rect 130 43697 1580 43727
rect 130 43611 1580 43641
rect 130 43525 1580 43555
rect 130 43439 1580 43469
rect 130 43353 1580 43383
rect 130 43267 1580 43297
rect 130 43181 1580 43211
rect 130 43095 1580 43125
rect 130 43009 1580 43039
rect 130 42923 1580 42953
rect 130 42837 1580 42867
rect 130 42751 1580 42781
rect 130 42665 1580 42695
rect 130 42579 1580 42609
rect 130 42493 1580 42523
rect 130 42407 1580 42437
rect 130 42321 1580 42351
rect 130 42235 1580 42265
rect 130 42149 1580 42179
rect 130 42063 1580 42093
rect 130 41977 1580 42007
rect 130 41891 1580 41921
rect 130 41805 1580 41835
rect 130 41719 1580 41749
rect 130 41633 1580 41663
rect 130 41547 1580 41577
rect 130 41461 1580 41491
rect 130 41375 1580 41405
rect 130 41289 1580 41319
rect 130 41203 1580 41233
rect 130 41117 1580 41147
rect 130 41031 1580 41061
rect 130 40945 1580 40975
rect 130 40859 1580 40889
rect 130 40773 1580 40803
rect 130 40687 1580 40717
rect 130 40601 1580 40631
rect 130 40515 1580 40545
rect 130 40429 1580 40459
rect 130 40343 1580 40373
rect 130 40257 1580 40287
rect 130 40171 1580 40201
rect 130 40085 1580 40115
rect 130 39999 1580 40029
rect 130 39913 1580 39943
rect 130 39827 1580 39857
rect 130 39741 1580 39771
rect 130 39655 1580 39685
rect 130 39569 1580 39599
rect 130 39483 1580 39513
rect 130 39397 1580 39427
rect 130 39311 1580 39341
rect 130 39225 1580 39255
rect 130 39139 1580 39169
rect 130 39053 1580 39083
rect 130 38967 1580 38997
rect 130 38881 1580 38911
rect 130 38795 1580 38825
rect 130 38709 1580 38739
rect 130 38623 1580 38653
rect 130 38537 1580 38567
rect 130 38451 1580 38481
rect 130 38365 1580 38395
rect 130 38279 1580 38309
rect 130 38193 1580 38223
rect 130 38107 1580 38137
rect 130 38021 1580 38051
rect 130 37935 1580 37965
rect 130 37849 1580 37879
rect 130 37763 1580 37793
rect 130 37677 1580 37707
rect 130 37591 1580 37621
rect 130 37505 1580 37535
rect 130 37419 1580 37449
rect 130 37333 1580 37363
rect 130 37247 1580 37277
rect 130 37161 1580 37191
rect 130 37075 1580 37105
rect 130 36989 1580 37019
rect 130 36903 1580 36933
rect 130 36817 1580 36847
rect 130 36731 1580 36761
rect 130 36645 1580 36675
rect 130 36559 1580 36589
rect 130 36473 1580 36503
rect 130 36387 1580 36417
rect 130 36301 1580 36331
rect 130 36215 1580 36245
rect 130 36129 1580 36159
rect 130 36043 1580 36073
rect 130 35957 1580 35987
rect 130 35871 1580 35901
rect 130 35785 1580 35815
rect 130 35699 1580 35729
rect 130 35613 1580 35643
rect 130 35527 1580 35557
rect 130 35441 1580 35471
rect 130 35355 1580 35385
rect 130 35269 1580 35299
rect 130 35183 1580 35213
rect 130 35097 1580 35127
rect 130 35011 1580 35041
rect 130 34925 1580 34955
rect 130 34839 1580 34869
rect 130 34753 1580 34783
rect 130 34667 1580 34697
rect 130 34581 1580 34611
rect 130 34495 1580 34525
rect 130 34409 1580 34439
rect 130 34323 1580 34353
rect 130 34237 1580 34267
rect 130 34151 1580 34181
rect 130 34065 1580 34095
rect 130 33979 1580 34009
rect 130 33893 1580 33923
rect 130 33807 1580 33837
rect 130 33721 1580 33751
rect 130 33635 1580 33665
rect 130 33549 1580 33579
rect 130 33463 1580 33493
rect 130 33377 1580 33407
rect 130 33291 1580 33321
rect 130 33205 1580 33235
rect 130 33119 1580 33149
rect 130 33033 1580 33063
rect 130 32947 1580 32977
rect 130 32861 1580 32891
rect 130 32775 1580 32805
rect 130 32689 1580 32719
rect 130 32603 1580 32633
rect 130 32517 1580 32547
rect 130 32431 1580 32461
rect 130 32345 1580 32375
rect 130 32259 1580 32289
rect 130 32173 1580 32203
rect 130 32087 1580 32117
rect 130 32001 1580 32031
rect 130 31915 1580 31945
rect 130 31829 1580 31859
rect 130 31743 1580 31773
rect 130 31657 1580 31687
rect 130 31571 1580 31601
rect 130 31485 1580 31515
rect 130 31399 1580 31429
rect 130 31313 1580 31343
rect 130 31227 1580 31257
rect 130 31141 1580 31171
rect 130 31055 1580 31085
rect 130 30969 1580 30999
rect 130 30883 1580 30913
rect 130 30797 1580 30827
rect 130 30711 1580 30741
rect 130 30625 1580 30655
rect 130 30539 1580 30569
rect 130 30453 1580 30483
rect 130 30367 1580 30397
rect 130 30281 1580 30311
rect 130 30195 1580 30225
rect 130 30109 1580 30139
rect 130 30023 1580 30053
rect 130 29937 1580 29967
rect 130 29851 1580 29881
rect 130 29765 1580 29795
rect 130 29679 1580 29709
rect 130 29593 1580 29623
rect 130 29507 1580 29537
rect 130 29421 1580 29451
rect 130 29335 1580 29365
rect 130 29249 1580 29279
rect 130 29163 1580 29193
rect 130 29077 1580 29107
rect 130 28991 1580 29021
rect 130 28905 1580 28935
rect 130 28819 1580 28849
rect 130 28733 1580 28763
rect 130 28647 1580 28677
rect 130 28561 1580 28591
rect 130 28475 1580 28505
rect 130 28389 1580 28419
rect 130 28303 1580 28333
rect 130 28217 1580 28247
rect 130 28131 1580 28161
rect 130 28045 1580 28075
rect 130 27959 1580 27989
rect 130 27873 1580 27903
rect 130 27787 1580 27817
rect 130 27701 1580 27731
rect 130 27615 1580 27645
rect 130 27529 1580 27559
rect 130 27443 1580 27473
rect 130 27357 1580 27387
rect 130 27271 1580 27301
rect 130 27185 1580 27215
rect 130 27099 1580 27129
rect 130 27013 1580 27043
rect 130 26927 1580 26957
rect 130 26841 1580 26871
rect 130 26755 1580 26785
rect 130 26669 1580 26699
rect 130 26583 1580 26613
rect 130 26497 1580 26527
rect 130 26411 1580 26441
rect 130 26325 1580 26355
rect 130 26239 1580 26269
rect 130 26153 1580 26183
rect 130 26067 1580 26097
rect 130 25981 1580 26011
rect 130 25895 1580 25925
rect 130 25809 1580 25839
rect 130 25723 1580 25753
rect 130 25637 1580 25667
rect 130 25551 1580 25581
rect 130 25465 1580 25495
rect 130 25379 1580 25409
rect 130 25293 1580 25323
rect 130 25207 1580 25237
rect 130 25121 1580 25151
rect 130 25035 1580 25065
rect 130 24949 1580 24979
rect 130 24863 1580 24893
rect 130 24777 1580 24807
rect 130 24691 1580 24721
rect 130 24605 1580 24635
rect 130 24519 1580 24549
rect 130 24433 1580 24463
rect 130 24347 1580 24377
rect 130 24261 1580 24291
rect 130 24175 1580 24205
rect 130 24089 1580 24119
rect 130 24003 1580 24033
rect 130 23917 1580 23947
rect 130 23831 1580 23861
rect 130 23745 1580 23775
rect 130 23659 1580 23689
rect 130 23573 1580 23603
rect 130 23487 1580 23517
rect 130 23401 1580 23431
rect 130 23315 1580 23345
rect 130 23229 1580 23259
rect 130 23143 1580 23173
rect 130 23057 1580 23087
rect 130 22971 1580 23001
rect 130 22885 1580 22915
rect 130 22799 1580 22829
rect 130 22713 1580 22743
rect 130 22627 1580 22657
rect 130 22541 1580 22571
rect 130 22455 1580 22485
rect 130 22369 1580 22399
rect 130 22283 1580 22313
rect 130 22197 1580 22227
rect 130 22111 1580 22141
rect 130 22025 1580 22055
rect 130 21939 1580 21969
rect 130 21853 1580 21883
rect 130 21767 1580 21797
rect 130 21681 1580 21711
rect 130 21595 1580 21625
rect 130 21509 1580 21539
rect 130 21423 1580 21453
rect 130 21337 1580 21367
rect 130 21251 1580 21281
rect 130 21165 1580 21195
rect 130 21079 1580 21109
rect 130 20993 1580 21023
rect 130 20907 1580 20937
rect 130 20821 1580 20851
rect 130 20735 1580 20765
rect 130 20649 1580 20679
rect 130 20563 1580 20593
rect 130 20477 1580 20507
rect 130 20391 1580 20421
rect 130 20305 1580 20335
rect 130 20219 1580 20249
rect 130 20133 1580 20163
rect 130 20047 1580 20077
rect 130 19961 1580 19991
rect 130 19875 1580 19905
rect 130 19789 1580 19819
rect 130 19703 1580 19733
rect 130 19617 1580 19647
rect 130 19531 1580 19561
rect 130 19445 1580 19475
rect 130 19359 1580 19389
rect 130 19273 1580 19303
rect 130 19187 1580 19217
rect 130 19101 1580 19131
rect 130 19015 1580 19045
rect 130 18929 1580 18959
rect 130 18843 1580 18873
rect 130 18757 1580 18787
rect 130 18671 1580 18701
rect 130 18585 1580 18615
rect 130 18499 1580 18529
rect 130 18413 1580 18443
rect 130 18327 1580 18357
rect 130 18241 1580 18271
rect 130 18155 1580 18185
rect 130 18069 1580 18099
rect 130 17983 1580 18013
rect 130 17897 1580 17927
rect 130 17811 1580 17841
rect 130 17725 1580 17755
rect 130 17639 1580 17669
rect 130 17553 1580 17583
rect 130 17467 1580 17497
rect 130 17381 1580 17411
rect 130 17295 1580 17325
rect 130 17209 1580 17239
rect 130 17123 1580 17153
rect 130 17037 1580 17067
rect 130 16951 1580 16981
rect 130 16865 1580 16895
rect 130 16779 1580 16809
rect 130 16693 1580 16723
rect 130 16607 1580 16637
rect 130 16521 1580 16551
rect 130 16435 1580 16465
rect 130 16349 1580 16379
rect 130 16263 1580 16293
rect 130 16177 1580 16207
rect 130 16091 1580 16121
rect 130 16005 1580 16035
rect 130 15919 1580 15949
rect 130 15833 1580 15863
rect 130 15747 1580 15777
rect 130 15661 1580 15691
rect 130 15575 1580 15605
rect 130 15489 1580 15519
rect 130 15403 1580 15433
rect 130 15317 1580 15347
rect 130 15231 1580 15261
rect 130 15145 1580 15175
rect 130 15059 1580 15089
rect 130 14973 1580 15003
rect 130 14887 1580 14917
rect 130 14801 1580 14831
rect 130 14715 1580 14745
rect 130 14629 1580 14659
rect 130 14543 1580 14573
rect 130 14457 1580 14487
rect 130 14371 1580 14401
rect 130 14285 1580 14315
rect 130 14199 1580 14229
rect 130 14113 1580 14143
rect 130 14027 1580 14057
rect 130 13941 1580 13971
rect 130 13855 1580 13885
rect 130 13769 1580 13799
rect 130 13683 1580 13713
rect 130 13597 1580 13627
rect 130 13511 1580 13541
rect 130 13425 1580 13455
rect 130 13339 1580 13369
rect 130 13253 1580 13283
rect 130 13167 1580 13197
rect 130 13081 1580 13111
rect 130 12995 1580 13025
rect 130 12909 1580 12939
rect 130 12823 1580 12853
rect 130 12737 1580 12767
rect 130 12651 1580 12681
rect 130 12565 1580 12595
rect 130 12479 1580 12509
rect 130 12393 1580 12423
rect 130 12307 1580 12337
rect 130 12221 1580 12251
rect 130 12135 1580 12165
rect 130 12049 1580 12079
rect 130 11963 1580 11993
rect 130 11877 1580 11907
rect 130 11791 1580 11821
rect 130 11705 1580 11735
rect 130 11619 1580 11649
rect 130 11533 1580 11563
rect 130 11447 1580 11477
rect 130 11361 1580 11391
rect 130 11275 1580 11305
rect 130 11189 1580 11219
rect 130 11103 1580 11133
rect 130 11017 1580 11047
rect 130 10931 1580 10961
rect 130 10845 1580 10875
rect 130 10759 1580 10789
rect 130 10673 1580 10703
rect 130 10587 1580 10617
rect 130 10501 1580 10531
rect 130 10415 1580 10445
rect 130 10329 1580 10359
rect 130 10243 1580 10273
rect 130 10157 1580 10187
rect 130 10071 1580 10101
rect 130 9985 1580 10015
rect 130 9899 1580 9929
rect 130 9813 1580 9843
rect 130 9727 1580 9757
rect 130 9641 1580 9671
rect 130 9555 1580 9585
rect 130 9469 1580 9499
rect 130 9383 1580 9413
rect 130 9297 1580 9327
rect 130 9211 1580 9241
rect 130 9125 1580 9155
rect 130 9039 1580 9069
rect 130 8953 1580 8983
rect 130 8867 1580 8897
rect 130 8781 1580 8811
rect 130 8695 1580 8725
rect 130 8609 1580 8639
rect 130 8523 1580 8553
rect 130 8437 1580 8467
rect 130 8351 1580 8381
rect 130 8265 1580 8295
rect 130 8179 1580 8209
rect 130 8093 1580 8123
rect 130 8007 1580 8037
rect 130 7921 1580 7951
rect 130 7835 1580 7865
rect 130 7749 1580 7779
rect 130 7663 1580 7693
rect 130 7577 1580 7607
rect 130 7491 1580 7521
rect 130 7405 1580 7435
rect 130 7319 1580 7349
rect 130 7233 1580 7263
rect 130 7147 1580 7177
rect 130 7061 1580 7091
rect 130 6975 1580 7005
rect 130 6889 1580 6919
rect 130 6803 1580 6833
rect 130 6717 1580 6747
rect 130 6631 1580 6661
rect 130 6545 1580 6575
rect 130 6459 1580 6489
rect 130 6373 1580 6403
rect 130 6287 1580 6317
rect 130 6201 1580 6231
rect 130 6115 1580 6145
rect 130 6029 1580 6059
rect 130 5943 1580 5973
rect 130 5857 1580 5887
rect 130 5771 1580 5801
rect 130 5685 1580 5715
rect 130 5599 1580 5629
rect 130 5513 1580 5543
rect 130 5427 1580 5457
rect 130 5341 1580 5371
rect 130 5255 1580 5285
rect 130 5169 1580 5199
rect 130 5083 1580 5113
rect 130 4997 1580 5027
rect 130 4911 1580 4941
rect 130 4825 1580 4855
rect 130 4739 1580 4769
rect 130 4653 1580 4683
rect 130 4567 1580 4597
rect 130 4481 1580 4511
rect 130 4395 1580 4425
rect 130 4309 1580 4339
rect 130 4223 1580 4253
rect 130 4137 1580 4167
rect 130 4051 1580 4081
rect 130 3965 1580 3995
rect 130 3879 1580 3909
rect 130 3793 1580 3823
rect 130 3707 1580 3737
rect 130 3621 1580 3651
rect 130 3535 1580 3565
rect 130 3449 1580 3479
rect 130 3363 1580 3393
rect 130 3277 1580 3307
rect 130 3191 1580 3221
rect 130 3105 1580 3135
rect 130 3019 1580 3049
rect 130 2933 1580 2963
rect 130 2847 1580 2877
rect 130 2761 1580 2791
rect 130 2675 1580 2705
rect 130 2589 1580 2619
rect 130 2503 1580 2533
rect 130 2417 1580 2447
rect 130 2331 1580 2361
rect 130 2245 1580 2275
rect 130 2159 1580 2189
rect 130 2073 1580 2103
rect 130 1987 1580 2017
rect 130 1901 1580 1931
rect 130 1815 1580 1845
rect 130 1729 1580 1759
rect 130 1643 1580 1673
rect 130 1557 1580 1587
rect 130 1471 1580 1501
rect 130 1385 1580 1415
rect 130 1299 1580 1329
rect 130 1213 1580 1243
rect 130 1127 1580 1157
rect 130 1041 1580 1071
rect 130 955 1580 985
rect 130 869 1580 899
rect 130 783 1580 813
rect 130 697 1580 727
rect 130 611 1580 641
rect 130 525 1580 555
rect 130 439 1580 469
rect 130 353 1580 383
rect 130 267 1580 297
rect 130 181 1580 211
<< pdiff >>
rect 130 100102 1580 100114
rect 130 100068 138 100102
rect 1572 100068 1580 100102
rect 130 100057 1580 100068
rect 130 100016 1580 100027
rect 130 99982 138 100016
rect 1572 99982 1580 100016
rect 130 99971 1580 99982
rect 130 99930 1580 99941
rect 130 99896 138 99930
rect 1572 99896 1580 99930
rect 130 99885 1580 99896
rect 130 99844 1580 99855
rect 130 99810 138 99844
rect 1572 99810 1580 99844
rect 130 99799 1580 99810
rect 130 99758 1580 99769
rect 130 99724 138 99758
rect 1572 99724 1580 99758
rect 130 99713 1580 99724
rect 130 99672 1580 99683
rect 130 99638 138 99672
rect 1572 99638 1580 99672
rect 130 99627 1580 99638
rect 130 99586 1580 99597
rect 130 99552 138 99586
rect 1572 99552 1580 99586
rect 130 99541 1580 99552
rect 130 99500 1580 99511
rect 130 99466 138 99500
rect 1572 99466 1580 99500
rect 130 99455 1580 99466
rect 130 99414 1580 99425
rect 130 99380 138 99414
rect 1572 99380 1580 99414
rect 130 99369 1580 99380
rect 130 99328 1580 99339
rect 130 99294 138 99328
rect 1572 99294 1580 99328
rect 130 99283 1580 99294
rect 130 99242 1580 99253
rect 130 99208 138 99242
rect 1572 99208 1580 99242
rect 130 99197 1580 99208
rect 130 99156 1580 99167
rect 130 99122 138 99156
rect 1572 99122 1580 99156
rect 130 99111 1580 99122
rect 130 99070 1580 99081
rect 130 99036 138 99070
rect 1572 99036 1580 99070
rect 130 99025 1580 99036
rect 130 98984 1580 98995
rect 130 98950 138 98984
rect 1572 98950 1580 98984
rect 130 98939 1580 98950
rect 130 98898 1580 98909
rect 130 98864 138 98898
rect 1572 98864 1580 98898
rect 130 98853 1580 98864
rect 130 98812 1580 98823
rect 130 98778 138 98812
rect 1572 98778 1580 98812
rect 130 98767 1580 98778
rect 130 98726 1580 98737
rect 130 98692 138 98726
rect 1572 98692 1580 98726
rect 130 98681 1580 98692
rect 130 98640 1580 98651
rect 130 98606 138 98640
rect 1572 98606 1580 98640
rect 130 98595 1580 98606
rect 130 98554 1580 98565
rect 130 98520 138 98554
rect 1572 98520 1580 98554
rect 130 98509 1580 98520
rect 130 98468 1580 98479
rect 130 98434 138 98468
rect 1572 98434 1580 98468
rect 130 98423 1580 98434
rect 130 98382 1580 98393
rect 130 98348 138 98382
rect 1572 98348 1580 98382
rect 130 98337 1580 98348
rect 130 98296 1580 98307
rect 130 98262 138 98296
rect 1572 98262 1580 98296
rect 130 98251 1580 98262
rect 130 98210 1580 98221
rect 130 98176 138 98210
rect 1572 98176 1580 98210
rect 130 98165 1580 98176
rect 130 98124 1580 98135
rect 130 98090 138 98124
rect 1572 98090 1580 98124
rect 130 98079 1580 98090
rect 130 98038 1580 98049
rect 130 98004 138 98038
rect 1572 98004 1580 98038
rect 130 97993 1580 98004
rect 130 97952 1580 97963
rect 130 97918 138 97952
rect 1572 97918 1580 97952
rect 130 97907 1580 97918
rect 130 97866 1580 97877
rect 130 97832 138 97866
rect 1572 97832 1580 97866
rect 130 97821 1580 97832
rect 130 97780 1580 97791
rect 130 97746 138 97780
rect 1572 97746 1580 97780
rect 130 97735 1580 97746
rect 130 97694 1580 97705
rect 130 97660 138 97694
rect 1572 97660 1580 97694
rect 130 97649 1580 97660
rect 130 97608 1580 97619
rect 130 97574 138 97608
rect 1572 97574 1580 97608
rect 130 97563 1580 97574
rect 130 97522 1580 97533
rect 130 97488 138 97522
rect 1572 97488 1580 97522
rect 130 97477 1580 97488
rect 130 97436 1580 97447
rect 130 97402 138 97436
rect 1572 97402 1580 97436
rect 130 97391 1580 97402
rect 130 97350 1580 97361
rect 130 97316 138 97350
rect 1572 97316 1580 97350
rect 130 97305 1580 97316
rect 130 97264 1580 97275
rect 130 97230 138 97264
rect 1572 97230 1580 97264
rect 130 97219 1580 97230
rect 130 97178 1580 97189
rect 130 97144 138 97178
rect 1572 97144 1580 97178
rect 130 97133 1580 97144
rect 130 97092 1580 97103
rect 130 97058 138 97092
rect 1572 97058 1580 97092
rect 130 97047 1580 97058
rect 130 97006 1580 97017
rect 130 96972 138 97006
rect 1572 96972 1580 97006
rect 130 96961 1580 96972
rect 130 96920 1580 96931
rect 130 96886 138 96920
rect 1572 96886 1580 96920
rect 130 96875 1580 96886
rect 130 96834 1580 96845
rect 130 96800 138 96834
rect 1572 96800 1580 96834
rect 130 96789 1580 96800
rect 130 96748 1580 96759
rect 130 96714 138 96748
rect 1572 96714 1580 96748
rect 130 96703 1580 96714
rect 130 96662 1580 96673
rect 130 96628 138 96662
rect 1572 96628 1580 96662
rect 130 96617 1580 96628
rect 130 96576 1580 96587
rect 130 96542 138 96576
rect 1572 96542 1580 96576
rect 130 96531 1580 96542
rect 130 96490 1580 96501
rect 130 96456 138 96490
rect 1572 96456 1580 96490
rect 130 96445 1580 96456
rect 130 96404 1580 96415
rect 130 96370 138 96404
rect 1572 96370 1580 96404
rect 130 96359 1580 96370
rect 130 96318 1580 96329
rect 130 96284 138 96318
rect 1572 96284 1580 96318
rect 130 96273 1580 96284
rect 130 96232 1580 96243
rect 130 96198 138 96232
rect 1572 96198 1580 96232
rect 130 96187 1580 96198
rect 130 96146 1580 96157
rect 130 96112 138 96146
rect 1572 96112 1580 96146
rect 130 96101 1580 96112
rect 130 96060 1580 96071
rect 130 96026 138 96060
rect 1572 96026 1580 96060
rect 130 96015 1580 96026
rect 130 95974 1580 95985
rect 130 95940 138 95974
rect 1572 95940 1580 95974
rect 130 95929 1580 95940
rect 130 95888 1580 95899
rect 130 95854 138 95888
rect 1572 95854 1580 95888
rect 130 95843 1580 95854
rect 130 95802 1580 95813
rect 130 95768 138 95802
rect 1572 95768 1580 95802
rect 130 95757 1580 95768
rect 130 95716 1580 95727
rect 130 95682 138 95716
rect 1572 95682 1580 95716
rect 130 95671 1580 95682
rect 130 95630 1580 95641
rect 130 95596 138 95630
rect 1572 95596 1580 95630
rect 130 95585 1580 95596
rect 130 95544 1580 95555
rect 130 95510 138 95544
rect 1572 95510 1580 95544
rect 130 95499 1580 95510
rect 130 95458 1580 95469
rect 130 95424 138 95458
rect 1572 95424 1580 95458
rect 130 95413 1580 95424
rect 130 95372 1580 95383
rect 130 95338 138 95372
rect 1572 95338 1580 95372
rect 130 95327 1580 95338
rect 130 95286 1580 95297
rect 130 95252 138 95286
rect 1572 95252 1580 95286
rect 130 95241 1580 95252
rect 130 95200 1580 95211
rect 130 95166 138 95200
rect 1572 95166 1580 95200
rect 130 95155 1580 95166
rect 130 95114 1580 95125
rect 130 95080 138 95114
rect 1572 95080 1580 95114
rect 130 95069 1580 95080
rect 130 95028 1580 95039
rect 130 94994 138 95028
rect 1572 94994 1580 95028
rect 130 94983 1580 94994
rect 130 94942 1580 94953
rect 130 94908 138 94942
rect 1572 94908 1580 94942
rect 130 94897 1580 94908
rect 130 94856 1580 94867
rect 130 94822 138 94856
rect 1572 94822 1580 94856
rect 130 94811 1580 94822
rect 130 94770 1580 94781
rect 130 94736 138 94770
rect 1572 94736 1580 94770
rect 130 94725 1580 94736
rect 130 94684 1580 94695
rect 130 94650 138 94684
rect 1572 94650 1580 94684
rect 130 94639 1580 94650
rect 130 94598 1580 94609
rect 130 94564 138 94598
rect 1572 94564 1580 94598
rect 130 94553 1580 94564
rect 130 94512 1580 94523
rect 130 94478 138 94512
rect 1572 94478 1580 94512
rect 130 94467 1580 94478
rect 130 94426 1580 94437
rect 130 94392 138 94426
rect 1572 94392 1580 94426
rect 130 94381 1580 94392
rect 130 94340 1580 94351
rect 130 94306 138 94340
rect 1572 94306 1580 94340
rect 130 94295 1580 94306
rect 130 94254 1580 94265
rect 130 94220 138 94254
rect 1572 94220 1580 94254
rect 130 94209 1580 94220
rect 130 94168 1580 94179
rect 130 94134 138 94168
rect 1572 94134 1580 94168
rect 130 94123 1580 94134
rect 130 94082 1580 94093
rect 130 94048 138 94082
rect 1572 94048 1580 94082
rect 130 94037 1580 94048
rect 130 93996 1580 94007
rect 130 93962 138 93996
rect 1572 93962 1580 93996
rect 130 93951 1580 93962
rect 130 93910 1580 93921
rect 130 93876 138 93910
rect 1572 93876 1580 93910
rect 130 93865 1580 93876
rect 130 93824 1580 93835
rect 130 93790 138 93824
rect 1572 93790 1580 93824
rect 130 93779 1580 93790
rect 130 93738 1580 93749
rect 130 93704 138 93738
rect 1572 93704 1580 93738
rect 130 93693 1580 93704
rect 130 93652 1580 93663
rect 130 93618 138 93652
rect 1572 93618 1580 93652
rect 130 93607 1580 93618
rect 130 93566 1580 93577
rect 130 93532 138 93566
rect 1572 93532 1580 93566
rect 130 93521 1580 93532
rect 130 93480 1580 93491
rect 130 93446 138 93480
rect 1572 93446 1580 93480
rect 130 93435 1580 93446
rect 130 93394 1580 93405
rect 130 93360 138 93394
rect 1572 93360 1580 93394
rect 130 93349 1580 93360
rect 130 93308 1580 93319
rect 130 93274 138 93308
rect 1572 93274 1580 93308
rect 130 93263 1580 93274
rect 130 93222 1580 93233
rect 130 93188 138 93222
rect 1572 93188 1580 93222
rect 130 93177 1580 93188
rect 130 93136 1580 93147
rect 130 93102 138 93136
rect 1572 93102 1580 93136
rect 130 93091 1580 93102
rect 130 93050 1580 93061
rect 130 93016 138 93050
rect 1572 93016 1580 93050
rect 130 93005 1580 93016
rect 130 92964 1580 92975
rect 130 92930 138 92964
rect 1572 92930 1580 92964
rect 130 92919 1580 92930
rect 130 92878 1580 92889
rect 130 92844 138 92878
rect 1572 92844 1580 92878
rect 130 92833 1580 92844
rect 130 92792 1580 92803
rect 130 92758 138 92792
rect 1572 92758 1580 92792
rect 130 92747 1580 92758
rect 130 92706 1580 92717
rect 130 92672 138 92706
rect 1572 92672 1580 92706
rect 130 92661 1580 92672
rect 130 92620 1580 92631
rect 130 92586 138 92620
rect 1572 92586 1580 92620
rect 130 92575 1580 92586
rect 130 92534 1580 92545
rect 130 92500 138 92534
rect 1572 92500 1580 92534
rect 130 92489 1580 92500
rect 130 92448 1580 92459
rect 130 92414 138 92448
rect 1572 92414 1580 92448
rect 130 92403 1580 92414
rect 130 92362 1580 92373
rect 130 92328 138 92362
rect 1572 92328 1580 92362
rect 130 92317 1580 92328
rect 130 92276 1580 92287
rect 130 92242 138 92276
rect 1572 92242 1580 92276
rect 130 92231 1580 92242
rect 130 92190 1580 92201
rect 130 92156 138 92190
rect 1572 92156 1580 92190
rect 130 92145 1580 92156
rect 130 92104 1580 92115
rect 130 92070 138 92104
rect 1572 92070 1580 92104
rect 130 92059 1580 92070
rect 130 92018 1580 92029
rect 130 91984 138 92018
rect 1572 91984 1580 92018
rect 130 91973 1580 91984
rect 130 91932 1580 91943
rect 130 91898 138 91932
rect 1572 91898 1580 91932
rect 130 91887 1580 91898
rect 130 91846 1580 91857
rect 130 91812 138 91846
rect 1572 91812 1580 91846
rect 130 91801 1580 91812
rect 130 91760 1580 91771
rect 130 91726 138 91760
rect 1572 91726 1580 91760
rect 130 91715 1580 91726
rect 130 91674 1580 91685
rect 130 91640 138 91674
rect 1572 91640 1580 91674
rect 130 91629 1580 91640
rect 130 91588 1580 91599
rect 130 91554 138 91588
rect 1572 91554 1580 91588
rect 130 91543 1580 91554
rect 130 91502 1580 91513
rect 130 91468 138 91502
rect 1572 91468 1580 91502
rect 130 91457 1580 91468
rect 130 91416 1580 91427
rect 130 91382 138 91416
rect 1572 91382 1580 91416
rect 130 91371 1580 91382
rect 130 91330 1580 91341
rect 130 91296 138 91330
rect 1572 91296 1580 91330
rect 130 91285 1580 91296
rect 130 91244 1580 91255
rect 130 91210 138 91244
rect 1572 91210 1580 91244
rect 130 91199 1580 91210
rect 130 91158 1580 91169
rect 130 91124 138 91158
rect 1572 91124 1580 91158
rect 130 91113 1580 91124
rect 130 91072 1580 91083
rect 130 91038 138 91072
rect 1572 91038 1580 91072
rect 130 91027 1580 91038
rect 130 90986 1580 90997
rect 130 90952 138 90986
rect 1572 90952 1580 90986
rect 130 90941 1580 90952
rect 130 90900 1580 90911
rect 130 90866 138 90900
rect 1572 90866 1580 90900
rect 130 90855 1580 90866
rect 130 90814 1580 90825
rect 130 90780 138 90814
rect 1572 90780 1580 90814
rect 130 90769 1580 90780
rect 130 90728 1580 90739
rect 130 90694 138 90728
rect 1572 90694 1580 90728
rect 130 90683 1580 90694
rect 130 90642 1580 90653
rect 130 90608 138 90642
rect 1572 90608 1580 90642
rect 130 90597 1580 90608
rect 130 90556 1580 90567
rect 130 90522 138 90556
rect 1572 90522 1580 90556
rect 130 90511 1580 90522
rect 130 90470 1580 90481
rect 130 90436 138 90470
rect 1572 90436 1580 90470
rect 130 90425 1580 90436
rect 130 90384 1580 90395
rect 130 90350 138 90384
rect 1572 90350 1580 90384
rect 130 90339 1580 90350
rect 130 90298 1580 90309
rect 130 90264 138 90298
rect 1572 90264 1580 90298
rect 130 90253 1580 90264
rect 130 90212 1580 90223
rect 130 90178 138 90212
rect 1572 90178 1580 90212
rect 130 90167 1580 90178
rect 130 90126 1580 90137
rect 130 90092 138 90126
rect 1572 90092 1580 90126
rect 130 90081 1580 90092
rect 130 90040 1580 90051
rect 130 90006 138 90040
rect 1572 90006 1580 90040
rect 130 89995 1580 90006
rect 130 89954 1580 89965
rect 130 89920 138 89954
rect 1572 89920 1580 89954
rect 130 89909 1580 89920
rect 130 89868 1580 89879
rect 130 89834 138 89868
rect 1572 89834 1580 89868
rect 130 89823 1580 89834
rect 130 89782 1580 89793
rect 130 89748 138 89782
rect 1572 89748 1580 89782
rect 130 89737 1580 89748
rect 130 89696 1580 89707
rect 130 89662 138 89696
rect 1572 89662 1580 89696
rect 130 89651 1580 89662
rect 130 89610 1580 89621
rect 130 89576 138 89610
rect 1572 89576 1580 89610
rect 130 89565 1580 89576
rect 130 89524 1580 89535
rect 130 89490 138 89524
rect 1572 89490 1580 89524
rect 130 89479 1580 89490
rect 130 89438 1580 89449
rect 130 89404 138 89438
rect 1572 89404 1580 89438
rect 130 89393 1580 89404
rect 130 89352 1580 89363
rect 130 89318 138 89352
rect 1572 89318 1580 89352
rect 130 89307 1580 89318
rect 130 89266 1580 89277
rect 130 89232 138 89266
rect 1572 89232 1580 89266
rect 130 89221 1580 89232
rect 130 89180 1580 89191
rect 130 89146 138 89180
rect 1572 89146 1580 89180
rect 130 89135 1580 89146
rect 130 89094 1580 89105
rect 130 89060 138 89094
rect 1572 89060 1580 89094
rect 130 89049 1580 89060
rect 130 89008 1580 89019
rect 130 88974 138 89008
rect 1572 88974 1580 89008
rect 130 88963 1580 88974
rect 130 88922 1580 88933
rect 130 88888 138 88922
rect 1572 88888 1580 88922
rect 130 88877 1580 88888
rect 130 88836 1580 88847
rect 130 88802 138 88836
rect 1572 88802 1580 88836
rect 130 88791 1580 88802
rect 130 88750 1580 88761
rect 130 88716 138 88750
rect 1572 88716 1580 88750
rect 130 88705 1580 88716
rect 130 88664 1580 88675
rect 130 88630 138 88664
rect 1572 88630 1580 88664
rect 130 88619 1580 88630
rect 130 88578 1580 88589
rect 130 88544 138 88578
rect 1572 88544 1580 88578
rect 130 88533 1580 88544
rect 130 88492 1580 88503
rect 130 88458 138 88492
rect 1572 88458 1580 88492
rect 130 88447 1580 88458
rect 130 88406 1580 88417
rect 130 88372 138 88406
rect 1572 88372 1580 88406
rect 130 88361 1580 88372
rect 130 88320 1580 88331
rect 130 88286 138 88320
rect 1572 88286 1580 88320
rect 130 88275 1580 88286
rect 130 88234 1580 88245
rect 130 88200 138 88234
rect 1572 88200 1580 88234
rect 130 88189 1580 88200
rect 130 88148 1580 88159
rect 130 88114 138 88148
rect 1572 88114 1580 88148
rect 130 88103 1580 88114
rect 130 88062 1580 88073
rect 130 88028 138 88062
rect 1572 88028 1580 88062
rect 130 88017 1580 88028
rect 130 87976 1580 87987
rect 130 87942 138 87976
rect 1572 87942 1580 87976
rect 130 87931 1580 87942
rect 130 87890 1580 87901
rect 130 87856 138 87890
rect 1572 87856 1580 87890
rect 130 87845 1580 87856
rect 130 87804 1580 87815
rect 130 87770 138 87804
rect 1572 87770 1580 87804
rect 130 87759 1580 87770
rect 130 87718 1580 87729
rect 130 87684 138 87718
rect 1572 87684 1580 87718
rect 130 87673 1580 87684
rect 130 87632 1580 87643
rect 130 87598 138 87632
rect 1572 87598 1580 87632
rect 130 87587 1580 87598
rect 130 87546 1580 87557
rect 130 87512 138 87546
rect 1572 87512 1580 87546
rect 130 87501 1580 87512
rect 130 87460 1580 87471
rect 130 87426 138 87460
rect 1572 87426 1580 87460
rect 130 87415 1580 87426
rect 130 87374 1580 87385
rect 130 87340 138 87374
rect 1572 87340 1580 87374
rect 130 87329 1580 87340
rect 130 87288 1580 87299
rect 130 87254 138 87288
rect 1572 87254 1580 87288
rect 130 87243 1580 87254
rect 130 87202 1580 87213
rect 130 87168 138 87202
rect 1572 87168 1580 87202
rect 130 87157 1580 87168
rect 130 87116 1580 87127
rect 130 87082 138 87116
rect 1572 87082 1580 87116
rect 130 87071 1580 87082
rect 130 87030 1580 87041
rect 130 86996 138 87030
rect 1572 86996 1580 87030
rect 130 86985 1580 86996
rect 130 86944 1580 86955
rect 130 86910 138 86944
rect 1572 86910 1580 86944
rect 130 86899 1580 86910
rect 130 86858 1580 86869
rect 130 86824 138 86858
rect 1572 86824 1580 86858
rect 130 86813 1580 86824
rect 130 86772 1580 86783
rect 130 86738 138 86772
rect 1572 86738 1580 86772
rect 130 86727 1580 86738
rect 130 86686 1580 86697
rect 130 86652 138 86686
rect 1572 86652 1580 86686
rect 130 86641 1580 86652
rect 130 86600 1580 86611
rect 130 86566 138 86600
rect 1572 86566 1580 86600
rect 130 86555 1580 86566
rect 130 86514 1580 86525
rect 130 86480 138 86514
rect 1572 86480 1580 86514
rect 130 86469 1580 86480
rect 130 86428 1580 86439
rect 130 86394 138 86428
rect 1572 86394 1580 86428
rect 130 86383 1580 86394
rect 130 86342 1580 86353
rect 130 86308 138 86342
rect 1572 86308 1580 86342
rect 130 86297 1580 86308
rect 130 86256 1580 86267
rect 130 86222 138 86256
rect 1572 86222 1580 86256
rect 130 86211 1580 86222
rect 130 86170 1580 86181
rect 130 86136 138 86170
rect 1572 86136 1580 86170
rect 130 86125 1580 86136
rect 130 86084 1580 86095
rect 130 86050 138 86084
rect 1572 86050 1580 86084
rect 130 86039 1580 86050
rect 130 85998 1580 86009
rect 130 85964 138 85998
rect 1572 85964 1580 85998
rect 130 85953 1580 85964
rect 130 85912 1580 85923
rect 130 85878 138 85912
rect 1572 85878 1580 85912
rect 130 85867 1580 85878
rect 130 85826 1580 85837
rect 130 85792 138 85826
rect 1572 85792 1580 85826
rect 130 85781 1580 85792
rect 130 85740 1580 85751
rect 130 85706 138 85740
rect 1572 85706 1580 85740
rect 130 85695 1580 85706
rect 130 85654 1580 85665
rect 130 85620 138 85654
rect 1572 85620 1580 85654
rect 130 85609 1580 85620
rect 130 85568 1580 85579
rect 130 85534 138 85568
rect 1572 85534 1580 85568
rect 130 85523 1580 85534
rect 130 85482 1580 85493
rect 130 85448 138 85482
rect 1572 85448 1580 85482
rect 130 85437 1580 85448
rect 130 85396 1580 85407
rect 130 85362 138 85396
rect 1572 85362 1580 85396
rect 130 85351 1580 85362
rect 130 85310 1580 85321
rect 130 85276 138 85310
rect 1572 85276 1580 85310
rect 130 85265 1580 85276
rect 130 85224 1580 85235
rect 130 85190 138 85224
rect 1572 85190 1580 85224
rect 130 85179 1580 85190
rect 130 85138 1580 85149
rect 130 85104 138 85138
rect 1572 85104 1580 85138
rect 130 85093 1580 85104
rect 130 85052 1580 85063
rect 130 85018 138 85052
rect 1572 85018 1580 85052
rect 130 85007 1580 85018
rect 130 84966 1580 84977
rect 130 84932 138 84966
rect 1572 84932 1580 84966
rect 130 84921 1580 84932
rect 130 84880 1580 84891
rect 130 84846 138 84880
rect 1572 84846 1580 84880
rect 130 84835 1580 84846
rect 130 84794 1580 84805
rect 130 84760 138 84794
rect 1572 84760 1580 84794
rect 130 84749 1580 84760
rect 130 84708 1580 84719
rect 130 84674 138 84708
rect 1572 84674 1580 84708
rect 130 84663 1580 84674
rect 130 84622 1580 84633
rect 130 84588 138 84622
rect 1572 84588 1580 84622
rect 130 84577 1580 84588
rect 130 84536 1580 84547
rect 130 84502 138 84536
rect 1572 84502 1580 84536
rect 130 84491 1580 84502
rect 130 84450 1580 84461
rect 130 84416 138 84450
rect 1572 84416 1580 84450
rect 130 84405 1580 84416
rect 130 84364 1580 84375
rect 130 84330 138 84364
rect 1572 84330 1580 84364
rect 130 84319 1580 84330
rect 130 84278 1580 84289
rect 130 84244 138 84278
rect 1572 84244 1580 84278
rect 130 84233 1580 84244
rect 130 84192 1580 84203
rect 130 84158 138 84192
rect 1572 84158 1580 84192
rect 130 84147 1580 84158
rect 130 84106 1580 84117
rect 130 84072 138 84106
rect 1572 84072 1580 84106
rect 130 84061 1580 84072
rect 130 84020 1580 84031
rect 130 83986 138 84020
rect 1572 83986 1580 84020
rect 130 83975 1580 83986
rect 130 83934 1580 83945
rect 130 83900 138 83934
rect 1572 83900 1580 83934
rect 130 83889 1580 83900
rect 130 83848 1580 83859
rect 130 83814 138 83848
rect 1572 83814 1580 83848
rect 130 83803 1580 83814
rect 130 83762 1580 83773
rect 130 83728 138 83762
rect 1572 83728 1580 83762
rect 130 83717 1580 83728
rect 130 83676 1580 83687
rect 130 83642 138 83676
rect 1572 83642 1580 83676
rect 130 83631 1580 83642
rect 130 83590 1580 83601
rect 130 83556 138 83590
rect 1572 83556 1580 83590
rect 130 83545 1580 83556
rect 130 83504 1580 83515
rect 130 83470 138 83504
rect 1572 83470 1580 83504
rect 130 83459 1580 83470
rect 130 83418 1580 83429
rect 130 83384 138 83418
rect 1572 83384 1580 83418
rect 130 83373 1580 83384
rect 130 83332 1580 83343
rect 130 83298 138 83332
rect 1572 83298 1580 83332
rect 130 83287 1580 83298
rect 130 83246 1580 83257
rect 130 83212 138 83246
rect 1572 83212 1580 83246
rect 130 83201 1580 83212
rect 130 83160 1580 83171
rect 130 83126 138 83160
rect 1572 83126 1580 83160
rect 130 83115 1580 83126
rect 130 83074 1580 83085
rect 130 83040 138 83074
rect 1572 83040 1580 83074
rect 130 83029 1580 83040
rect 130 82988 1580 82999
rect 130 82954 138 82988
rect 1572 82954 1580 82988
rect 130 82943 1580 82954
rect 130 82902 1580 82913
rect 130 82868 138 82902
rect 1572 82868 1580 82902
rect 130 82857 1580 82868
rect 130 82816 1580 82827
rect 130 82782 138 82816
rect 1572 82782 1580 82816
rect 130 82771 1580 82782
rect 130 82730 1580 82741
rect 130 82696 138 82730
rect 1572 82696 1580 82730
rect 130 82685 1580 82696
rect 130 82644 1580 82655
rect 130 82610 138 82644
rect 1572 82610 1580 82644
rect 130 82599 1580 82610
rect 130 82558 1580 82569
rect 130 82524 138 82558
rect 1572 82524 1580 82558
rect 130 82513 1580 82524
rect 130 82472 1580 82483
rect 130 82438 138 82472
rect 1572 82438 1580 82472
rect 130 82427 1580 82438
rect 130 82386 1580 82397
rect 130 82352 138 82386
rect 1572 82352 1580 82386
rect 130 82341 1580 82352
rect 130 82300 1580 82311
rect 130 82266 138 82300
rect 1572 82266 1580 82300
rect 130 82255 1580 82266
rect 130 82214 1580 82225
rect 130 82180 138 82214
rect 1572 82180 1580 82214
rect 130 82169 1580 82180
rect 130 82128 1580 82139
rect 130 82094 138 82128
rect 1572 82094 1580 82128
rect 130 82083 1580 82094
rect 130 82042 1580 82053
rect 130 82008 138 82042
rect 1572 82008 1580 82042
rect 130 81997 1580 82008
rect 130 81956 1580 81967
rect 130 81922 138 81956
rect 1572 81922 1580 81956
rect 130 81911 1580 81922
rect 130 81870 1580 81881
rect 130 81836 138 81870
rect 1572 81836 1580 81870
rect 130 81825 1580 81836
rect 130 81784 1580 81795
rect 130 81750 138 81784
rect 1572 81750 1580 81784
rect 130 81739 1580 81750
rect 130 81698 1580 81709
rect 130 81664 138 81698
rect 1572 81664 1580 81698
rect 130 81653 1580 81664
rect 130 81612 1580 81623
rect 130 81578 138 81612
rect 1572 81578 1580 81612
rect 130 81567 1580 81578
rect 130 81526 1580 81537
rect 130 81492 138 81526
rect 1572 81492 1580 81526
rect 130 81481 1580 81492
rect 130 81440 1580 81451
rect 130 81406 138 81440
rect 1572 81406 1580 81440
rect 130 81395 1580 81406
rect 130 81354 1580 81365
rect 130 81320 138 81354
rect 1572 81320 1580 81354
rect 130 81309 1580 81320
rect 130 81268 1580 81279
rect 130 81234 138 81268
rect 1572 81234 1580 81268
rect 130 81223 1580 81234
rect 130 81182 1580 81193
rect 130 81148 138 81182
rect 1572 81148 1580 81182
rect 130 81137 1580 81148
rect 130 81096 1580 81107
rect 130 81062 138 81096
rect 1572 81062 1580 81096
rect 130 81051 1580 81062
rect 130 81010 1580 81021
rect 130 80976 138 81010
rect 1572 80976 1580 81010
rect 130 80965 1580 80976
rect 130 80924 1580 80935
rect 130 80890 138 80924
rect 1572 80890 1580 80924
rect 130 80879 1580 80890
rect 130 80838 1580 80849
rect 130 80804 138 80838
rect 1572 80804 1580 80838
rect 130 80793 1580 80804
rect 130 80752 1580 80763
rect 130 80718 138 80752
rect 1572 80718 1580 80752
rect 130 80707 1580 80718
rect 130 80666 1580 80677
rect 130 80632 138 80666
rect 1572 80632 1580 80666
rect 130 80621 1580 80632
rect 130 80580 1580 80591
rect 130 80546 138 80580
rect 1572 80546 1580 80580
rect 130 80535 1580 80546
rect 130 80494 1580 80505
rect 130 80460 138 80494
rect 1572 80460 1580 80494
rect 130 80449 1580 80460
rect 130 80408 1580 80419
rect 130 80374 138 80408
rect 1572 80374 1580 80408
rect 130 80363 1580 80374
rect 130 80322 1580 80333
rect 130 80288 138 80322
rect 1572 80288 1580 80322
rect 130 80277 1580 80288
rect 130 80236 1580 80247
rect 130 80202 138 80236
rect 1572 80202 1580 80236
rect 130 80191 1580 80202
rect 130 80150 1580 80161
rect 130 80116 138 80150
rect 1572 80116 1580 80150
rect 130 80105 1580 80116
rect 130 80064 1580 80075
rect 130 80030 138 80064
rect 1572 80030 1580 80064
rect 130 80019 1580 80030
rect 130 79978 1580 79989
rect 130 79944 138 79978
rect 1572 79944 1580 79978
rect 130 79933 1580 79944
rect 130 79892 1580 79903
rect 130 79858 138 79892
rect 1572 79858 1580 79892
rect 130 79847 1580 79858
rect 130 79806 1580 79817
rect 130 79772 138 79806
rect 1572 79772 1580 79806
rect 130 79761 1580 79772
rect 130 79720 1580 79731
rect 130 79686 138 79720
rect 1572 79686 1580 79720
rect 130 79675 1580 79686
rect 130 79634 1580 79645
rect 130 79600 138 79634
rect 1572 79600 1580 79634
rect 130 79589 1580 79600
rect 130 79548 1580 79559
rect 130 79514 138 79548
rect 1572 79514 1580 79548
rect 130 79503 1580 79514
rect 130 79462 1580 79473
rect 130 79428 138 79462
rect 1572 79428 1580 79462
rect 130 79417 1580 79428
rect 130 79376 1580 79387
rect 130 79342 138 79376
rect 1572 79342 1580 79376
rect 130 79331 1580 79342
rect 130 79290 1580 79301
rect 130 79256 138 79290
rect 1572 79256 1580 79290
rect 130 79245 1580 79256
rect 130 79204 1580 79215
rect 130 79170 138 79204
rect 1572 79170 1580 79204
rect 130 79159 1580 79170
rect 130 79118 1580 79129
rect 130 79084 138 79118
rect 1572 79084 1580 79118
rect 130 79073 1580 79084
rect 130 79032 1580 79043
rect 130 78998 138 79032
rect 1572 78998 1580 79032
rect 130 78987 1580 78998
rect 130 78946 1580 78957
rect 130 78912 138 78946
rect 1572 78912 1580 78946
rect 130 78901 1580 78912
rect 130 78860 1580 78871
rect 130 78826 138 78860
rect 1572 78826 1580 78860
rect 130 78815 1580 78826
rect 130 78774 1580 78785
rect 130 78740 138 78774
rect 1572 78740 1580 78774
rect 130 78729 1580 78740
rect 130 78688 1580 78699
rect 130 78654 138 78688
rect 1572 78654 1580 78688
rect 130 78643 1580 78654
rect 130 78602 1580 78613
rect 130 78568 138 78602
rect 1572 78568 1580 78602
rect 130 78557 1580 78568
rect 130 78516 1580 78527
rect 130 78482 138 78516
rect 1572 78482 1580 78516
rect 130 78471 1580 78482
rect 130 78430 1580 78441
rect 130 78396 138 78430
rect 1572 78396 1580 78430
rect 130 78385 1580 78396
rect 130 78344 1580 78355
rect 130 78310 138 78344
rect 1572 78310 1580 78344
rect 130 78299 1580 78310
rect 130 78258 1580 78269
rect 130 78224 138 78258
rect 1572 78224 1580 78258
rect 130 78213 1580 78224
rect 130 78172 1580 78183
rect 130 78138 138 78172
rect 1572 78138 1580 78172
rect 130 78127 1580 78138
rect 130 78086 1580 78097
rect 130 78052 138 78086
rect 1572 78052 1580 78086
rect 130 78041 1580 78052
rect 130 78000 1580 78011
rect 130 77966 138 78000
rect 1572 77966 1580 78000
rect 130 77955 1580 77966
rect 130 77914 1580 77925
rect 130 77880 138 77914
rect 1572 77880 1580 77914
rect 130 77869 1580 77880
rect 130 77828 1580 77839
rect 130 77794 138 77828
rect 1572 77794 1580 77828
rect 130 77783 1580 77794
rect 130 77742 1580 77753
rect 130 77708 138 77742
rect 1572 77708 1580 77742
rect 130 77697 1580 77708
rect 130 77656 1580 77667
rect 130 77622 138 77656
rect 1572 77622 1580 77656
rect 130 77611 1580 77622
rect 130 77570 1580 77581
rect 130 77536 138 77570
rect 1572 77536 1580 77570
rect 130 77525 1580 77536
rect 130 77484 1580 77495
rect 130 77450 138 77484
rect 1572 77450 1580 77484
rect 130 77439 1580 77450
rect 130 77398 1580 77409
rect 130 77364 138 77398
rect 1572 77364 1580 77398
rect 130 77353 1580 77364
rect 130 77312 1580 77323
rect 130 77278 138 77312
rect 1572 77278 1580 77312
rect 130 77267 1580 77278
rect 130 77226 1580 77237
rect 130 77192 138 77226
rect 1572 77192 1580 77226
rect 130 77181 1580 77192
rect 130 77140 1580 77151
rect 130 77106 138 77140
rect 1572 77106 1580 77140
rect 130 77095 1580 77106
rect 130 77054 1580 77065
rect 130 77020 138 77054
rect 1572 77020 1580 77054
rect 130 77009 1580 77020
rect 130 76968 1580 76979
rect 130 76934 138 76968
rect 1572 76934 1580 76968
rect 130 76923 1580 76934
rect 130 76882 1580 76893
rect 130 76848 138 76882
rect 1572 76848 1580 76882
rect 130 76837 1580 76848
rect 130 76796 1580 76807
rect 130 76762 138 76796
rect 1572 76762 1580 76796
rect 130 76751 1580 76762
rect 130 76710 1580 76721
rect 130 76676 138 76710
rect 1572 76676 1580 76710
rect 130 76665 1580 76676
rect 130 76624 1580 76635
rect 130 76590 138 76624
rect 1572 76590 1580 76624
rect 130 76579 1580 76590
rect 130 76538 1580 76549
rect 130 76504 138 76538
rect 1572 76504 1580 76538
rect 130 76493 1580 76504
rect 130 76452 1580 76463
rect 130 76418 138 76452
rect 1572 76418 1580 76452
rect 130 76407 1580 76418
rect 130 76366 1580 76377
rect 130 76332 138 76366
rect 1572 76332 1580 76366
rect 130 76321 1580 76332
rect 130 76280 1580 76291
rect 130 76246 138 76280
rect 1572 76246 1580 76280
rect 130 76235 1580 76246
rect 130 76194 1580 76205
rect 130 76160 138 76194
rect 1572 76160 1580 76194
rect 130 76149 1580 76160
rect 130 76108 1580 76119
rect 130 76074 138 76108
rect 1572 76074 1580 76108
rect 130 76063 1580 76074
rect 130 76022 1580 76033
rect 130 75988 138 76022
rect 1572 75988 1580 76022
rect 130 75977 1580 75988
rect 130 75936 1580 75947
rect 130 75902 138 75936
rect 1572 75902 1580 75936
rect 130 75891 1580 75902
rect 130 75850 1580 75861
rect 130 75816 138 75850
rect 1572 75816 1580 75850
rect 130 75805 1580 75816
rect 130 75764 1580 75775
rect 130 75730 138 75764
rect 1572 75730 1580 75764
rect 130 75719 1580 75730
rect 130 75678 1580 75689
rect 130 75644 138 75678
rect 1572 75644 1580 75678
rect 130 75633 1580 75644
rect 130 75592 1580 75603
rect 130 75558 138 75592
rect 1572 75558 1580 75592
rect 130 75547 1580 75558
rect 130 75506 1580 75517
rect 130 75472 138 75506
rect 1572 75472 1580 75506
rect 130 75461 1580 75472
rect 130 75420 1580 75431
rect 130 75386 138 75420
rect 1572 75386 1580 75420
rect 130 75375 1580 75386
rect 130 75334 1580 75345
rect 130 75300 138 75334
rect 1572 75300 1580 75334
rect 130 75289 1580 75300
rect 130 75248 1580 75259
rect 130 75214 138 75248
rect 1572 75214 1580 75248
rect 130 75203 1580 75214
rect 130 75162 1580 75173
rect 130 75128 138 75162
rect 1572 75128 1580 75162
rect 130 75117 1580 75128
rect 130 75076 1580 75087
rect 130 75042 138 75076
rect 1572 75042 1580 75076
rect 130 75031 1580 75042
rect 130 74990 1580 75001
rect 130 74956 138 74990
rect 1572 74956 1580 74990
rect 130 74945 1580 74956
rect 130 74904 1580 74915
rect 130 74870 138 74904
rect 1572 74870 1580 74904
rect 130 74859 1580 74870
rect 130 74818 1580 74829
rect 130 74784 138 74818
rect 1572 74784 1580 74818
rect 130 74773 1580 74784
rect 130 74732 1580 74743
rect 130 74698 138 74732
rect 1572 74698 1580 74732
rect 130 74687 1580 74698
rect 130 74646 1580 74657
rect 130 74612 138 74646
rect 1572 74612 1580 74646
rect 130 74601 1580 74612
rect 130 74560 1580 74571
rect 130 74526 138 74560
rect 1572 74526 1580 74560
rect 130 74515 1580 74526
rect 130 74474 1580 74485
rect 130 74440 138 74474
rect 1572 74440 1580 74474
rect 130 74429 1580 74440
rect 130 74388 1580 74399
rect 130 74354 138 74388
rect 1572 74354 1580 74388
rect 130 74343 1580 74354
rect 130 74302 1580 74313
rect 130 74268 138 74302
rect 1572 74268 1580 74302
rect 130 74257 1580 74268
rect 130 74216 1580 74227
rect 130 74182 138 74216
rect 1572 74182 1580 74216
rect 130 74171 1580 74182
rect 130 74130 1580 74141
rect 130 74096 138 74130
rect 1572 74096 1580 74130
rect 130 74085 1580 74096
rect 130 74044 1580 74055
rect 130 74010 138 74044
rect 1572 74010 1580 74044
rect 130 73999 1580 74010
rect 130 73958 1580 73969
rect 130 73924 138 73958
rect 1572 73924 1580 73958
rect 130 73913 1580 73924
rect 130 73872 1580 73883
rect 130 73838 138 73872
rect 1572 73838 1580 73872
rect 130 73827 1580 73838
rect 130 73786 1580 73797
rect 130 73752 138 73786
rect 1572 73752 1580 73786
rect 130 73741 1580 73752
rect 130 73700 1580 73711
rect 130 73666 138 73700
rect 1572 73666 1580 73700
rect 130 73655 1580 73666
rect 130 73614 1580 73625
rect 130 73580 138 73614
rect 1572 73580 1580 73614
rect 130 73569 1580 73580
rect 130 73528 1580 73539
rect 130 73494 138 73528
rect 1572 73494 1580 73528
rect 130 73483 1580 73494
rect 130 73442 1580 73453
rect 130 73408 138 73442
rect 1572 73408 1580 73442
rect 130 73397 1580 73408
rect 130 73356 1580 73367
rect 130 73322 138 73356
rect 1572 73322 1580 73356
rect 130 73311 1580 73322
rect 130 73270 1580 73281
rect 130 73236 138 73270
rect 1572 73236 1580 73270
rect 130 73225 1580 73236
rect 130 73184 1580 73195
rect 130 73150 138 73184
rect 1572 73150 1580 73184
rect 130 73139 1580 73150
rect 130 73098 1580 73109
rect 130 73064 138 73098
rect 1572 73064 1580 73098
rect 130 73053 1580 73064
rect 130 73012 1580 73023
rect 130 72978 138 73012
rect 1572 72978 1580 73012
rect 130 72967 1580 72978
rect 130 72926 1580 72937
rect 130 72892 138 72926
rect 1572 72892 1580 72926
rect 130 72881 1580 72892
rect 130 72840 1580 72851
rect 130 72806 138 72840
rect 1572 72806 1580 72840
rect 130 72795 1580 72806
rect 130 72754 1580 72765
rect 130 72720 138 72754
rect 1572 72720 1580 72754
rect 130 72709 1580 72720
rect 130 72668 1580 72679
rect 130 72634 138 72668
rect 1572 72634 1580 72668
rect 130 72623 1580 72634
rect 130 72582 1580 72593
rect 130 72548 138 72582
rect 1572 72548 1580 72582
rect 130 72537 1580 72548
rect 130 72496 1580 72507
rect 130 72462 138 72496
rect 1572 72462 1580 72496
rect 130 72451 1580 72462
rect 130 72410 1580 72421
rect 130 72376 138 72410
rect 1572 72376 1580 72410
rect 130 72365 1580 72376
rect 130 72324 1580 72335
rect 130 72290 138 72324
rect 1572 72290 1580 72324
rect 130 72279 1580 72290
rect 130 72238 1580 72249
rect 130 72204 138 72238
rect 1572 72204 1580 72238
rect 130 72193 1580 72204
rect 130 72152 1580 72163
rect 130 72118 138 72152
rect 1572 72118 1580 72152
rect 130 72107 1580 72118
rect 130 72066 1580 72077
rect 130 72032 138 72066
rect 1572 72032 1580 72066
rect 130 72021 1580 72032
rect 130 71980 1580 71991
rect 130 71946 138 71980
rect 1572 71946 1580 71980
rect 130 71935 1580 71946
rect 130 71894 1580 71905
rect 130 71860 138 71894
rect 1572 71860 1580 71894
rect 130 71849 1580 71860
rect 130 71808 1580 71819
rect 130 71774 138 71808
rect 1572 71774 1580 71808
rect 130 71763 1580 71774
rect 130 71722 1580 71733
rect 130 71688 138 71722
rect 1572 71688 1580 71722
rect 130 71677 1580 71688
rect 130 71636 1580 71647
rect 130 71602 138 71636
rect 1572 71602 1580 71636
rect 130 71591 1580 71602
rect 130 71550 1580 71561
rect 130 71516 138 71550
rect 1572 71516 1580 71550
rect 130 71505 1580 71516
rect 130 71464 1580 71475
rect 130 71430 138 71464
rect 1572 71430 1580 71464
rect 130 71419 1580 71430
rect 130 71378 1580 71389
rect 130 71344 138 71378
rect 1572 71344 1580 71378
rect 130 71333 1580 71344
rect 130 71292 1580 71303
rect 130 71258 138 71292
rect 1572 71258 1580 71292
rect 130 71247 1580 71258
rect 130 71206 1580 71217
rect 130 71172 138 71206
rect 1572 71172 1580 71206
rect 130 71161 1580 71172
rect 130 71120 1580 71131
rect 130 71086 138 71120
rect 1572 71086 1580 71120
rect 130 71075 1580 71086
rect 130 71034 1580 71045
rect 130 71000 138 71034
rect 1572 71000 1580 71034
rect 130 70989 1580 71000
rect 130 70948 1580 70959
rect 130 70914 138 70948
rect 1572 70914 1580 70948
rect 130 70903 1580 70914
rect 130 70862 1580 70873
rect 130 70828 138 70862
rect 1572 70828 1580 70862
rect 130 70817 1580 70828
rect 130 70776 1580 70787
rect 130 70742 138 70776
rect 1572 70742 1580 70776
rect 130 70731 1580 70742
rect 130 70690 1580 70701
rect 130 70656 138 70690
rect 1572 70656 1580 70690
rect 130 70645 1580 70656
rect 130 70604 1580 70615
rect 130 70570 138 70604
rect 1572 70570 1580 70604
rect 130 70559 1580 70570
rect 130 70518 1580 70529
rect 130 70484 138 70518
rect 1572 70484 1580 70518
rect 130 70473 1580 70484
rect 130 70432 1580 70443
rect 130 70398 138 70432
rect 1572 70398 1580 70432
rect 130 70387 1580 70398
rect 130 70346 1580 70357
rect 130 70312 138 70346
rect 1572 70312 1580 70346
rect 130 70301 1580 70312
rect 130 70260 1580 70271
rect 130 70226 138 70260
rect 1572 70226 1580 70260
rect 130 70215 1580 70226
rect 130 70174 1580 70185
rect 130 70140 138 70174
rect 1572 70140 1580 70174
rect 130 70129 1580 70140
rect 130 70088 1580 70099
rect 130 70054 138 70088
rect 1572 70054 1580 70088
rect 130 70043 1580 70054
rect 130 70002 1580 70013
rect 130 69968 138 70002
rect 1572 69968 1580 70002
rect 130 69957 1580 69968
rect 130 69916 1580 69927
rect 130 69882 138 69916
rect 1572 69882 1580 69916
rect 130 69871 1580 69882
rect 130 69830 1580 69841
rect 130 69796 138 69830
rect 1572 69796 1580 69830
rect 130 69785 1580 69796
rect 130 69744 1580 69755
rect 130 69710 138 69744
rect 1572 69710 1580 69744
rect 130 69699 1580 69710
rect 130 69658 1580 69669
rect 130 69624 138 69658
rect 1572 69624 1580 69658
rect 130 69613 1580 69624
rect 130 69572 1580 69583
rect 130 69538 138 69572
rect 1572 69538 1580 69572
rect 130 69527 1580 69538
rect 130 69486 1580 69497
rect 130 69452 138 69486
rect 1572 69452 1580 69486
rect 130 69441 1580 69452
rect 130 69400 1580 69411
rect 130 69366 138 69400
rect 1572 69366 1580 69400
rect 130 69355 1580 69366
rect 130 69314 1580 69325
rect 130 69280 138 69314
rect 1572 69280 1580 69314
rect 130 69269 1580 69280
rect 130 69228 1580 69239
rect 130 69194 138 69228
rect 1572 69194 1580 69228
rect 130 69183 1580 69194
rect 130 69142 1580 69153
rect 130 69108 138 69142
rect 1572 69108 1580 69142
rect 130 69097 1580 69108
rect 130 69056 1580 69067
rect 130 69022 138 69056
rect 1572 69022 1580 69056
rect 130 69011 1580 69022
rect 130 68970 1580 68981
rect 130 68936 138 68970
rect 1572 68936 1580 68970
rect 130 68925 1580 68936
rect 130 68884 1580 68895
rect 130 68850 138 68884
rect 1572 68850 1580 68884
rect 130 68839 1580 68850
rect 130 68798 1580 68809
rect 130 68764 138 68798
rect 1572 68764 1580 68798
rect 130 68753 1580 68764
rect 130 68712 1580 68723
rect 130 68678 138 68712
rect 1572 68678 1580 68712
rect 130 68667 1580 68678
rect 130 68626 1580 68637
rect 130 68592 138 68626
rect 1572 68592 1580 68626
rect 130 68581 1580 68592
rect 130 68540 1580 68551
rect 130 68506 138 68540
rect 1572 68506 1580 68540
rect 130 68495 1580 68506
rect 130 68454 1580 68465
rect 130 68420 138 68454
rect 1572 68420 1580 68454
rect 130 68409 1580 68420
rect 130 68368 1580 68379
rect 130 68334 138 68368
rect 1572 68334 1580 68368
rect 130 68323 1580 68334
rect 130 68282 1580 68293
rect 130 68248 138 68282
rect 1572 68248 1580 68282
rect 130 68237 1580 68248
rect 130 68196 1580 68207
rect 130 68162 138 68196
rect 1572 68162 1580 68196
rect 130 68151 1580 68162
rect 130 68110 1580 68121
rect 130 68076 138 68110
rect 1572 68076 1580 68110
rect 130 68065 1580 68076
rect 130 68024 1580 68035
rect 130 67990 138 68024
rect 1572 67990 1580 68024
rect 130 67979 1580 67990
rect 130 67938 1580 67949
rect 130 67904 138 67938
rect 1572 67904 1580 67938
rect 130 67893 1580 67904
rect 130 67852 1580 67863
rect 130 67818 138 67852
rect 1572 67818 1580 67852
rect 130 67807 1580 67818
rect 130 67766 1580 67777
rect 130 67732 138 67766
rect 1572 67732 1580 67766
rect 130 67721 1580 67732
rect 130 67680 1580 67691
rect 130 67646 138 67680
rect 1572 67646 1580 67680
rect 130 67635 1580 67646
rect 130 67594 1580 67605
rect 130 67560 138 67594
rect 1572 67560 1580 67594
rect 130 67549 1580 67560
rect 130 67508 1580 67519
rect 130 67474 138 67508
rect 1572 67474 1580 67508
rect 130 67463 1580 67474
rect 130 67422 1580 67433
rect 130 67388 138 67422
rect 1572 67388 1580 67422
rect 130 67377 1580 67388
rect 130 67336 1580 67347
rect 130 67302 138 67336
rect 1572 67302 1580 67336
rect 130 67291 1580 67302
rect 130 67250 1580 67261
rect 130 67216 138 67250
rect 1572 67216 1580 67250
rect 130 67205 1580 67216
rect 130 67164 1580 67175
rect 130 67130 138 67164
rect 1572 67130 1580 67164
rect 130 67119 1580 67130
rect 130 67078 1580 67089
rect 130 67044 138 67078
rect 1572 67044 1580 67078
rect 130 67033 1580 67044
rect 130 66992 1580 67003
rect 130 66958 138 66992
rect 1572 66958 1580 66992
rect 130 66947 1580 66958
rect 130 66906 1580 66917
rect 130 66872 138 66906
rect 1572 66872 1580 66906
rect 130 66861 1580 66872
rect 130 66820 1580 66831
rect 130 66786 138 66820
rect 1572 66786 1580 66820
rect 130 66775 1580 66786
rect 130 66734 1580 66745
rect 130 66700 138 66734
rect 1572 66700 1580 66734
rect 130 66689 1580 66700
rect 130 66648 1580 66659
rect 130 66614 138 66648
rect 1572 66614 1580 66648
rect 130 66603 1580 66614
rect 130 66562 1580 66573
rect 130 66528 138 66562
rect 1572 66528 1580 66562
rect 130 66517 1580 66528
rect 130 66476 1580 66487
rect 130 66442 138 66476
rect 1572 66442 1580 66476
rect 130 66431 1580 66442
rect 130 66390 1580 66401
rect 130 66356 138 66390
rect 1572 66356 1580 66390
rect 130 66345 1580 66356
rect 130 66304 1580 66315
rect 130 66270 138 66304
rect 1572 66270 1580 66304
rect 130 66259 1580 66270
rect 130 66218 1580 66229
rect 130 66184 138 66218
rect 1572 66184 1580 66218
rect 130 66173 1580 66184
rect 130 66132 1580 66143
rect 130 66098 138 66132
rect 1572 66098 1580 66132
rect 130 66087 1580 66098
rect 130 66046 1580 66057
rect 130 66012 138 66046
rect 1572 66012 1580 66046
rect 130 66001 1580 66012
rect 130 65960 1580 65971
rect 130 65926 138 65960
rect 1572 65926 1580 65960
rect 130 65915 1580 65926
rect 130 65874 1580 65885
rect 130 65840 138 65874
rect 1572 65840 1580 65874
rect 130 65829 1580 65840
rect 130 65788 1580 65799
rect 130 65754 138 65788
rect 1572 65754 1580 65788
rect 130 65743 1580 65754
rect 130 65702 1580 65713
rect 130 65668 138 65702
rect 1572 65668 1580 65702
rect 130 65657 1580 65668
rect 130 65616 1580 65627
rect 130 65582 138 65616
rect 1572 65582 1580 65616
rect 130 65571 1580 65582
rect 130 65530 1580 65541
rect 130 65496 138 65530
rect 1572 65496 1580 65530
rect 130 65485 1580 65496
rect 130 65444 1580 65455
rect 130 65410 138 65444
rect 1572 65410 1580 65444
rect 130 65399 1580 65410
rect 130 65358 1580 65369
rect 130 65324 138 65358
rect 1572 65324 1580 65358
rect 130 65313 1580 65324
rect 130 65272 1580 65283
rect 130 65238 138 65272
rect 1572 65238 1580 65272
rect 130 65227 1580 65238
rect 130 65186 1580 65197
rect 130 65152 138 65186
rect 1572 65152 1580 65186
rect 130 65141 1580 65152
rect 130 65100 1580 65111
rect 130 65066 138 65100
rect 1572 65066 1580 65100
rect 130 65055 1580 65066
rect 130 65014 1580 65025
rect 130 64980 138 65014
rect 1572 64980 1580 65014
rect 130 64969 1580 64980
rect 130 64928 1580 64939
rect 130 64894 138 64928
rect 1572 64894 1580 64928
rect 130 64883 1580 64894
rect 130 64842 1580 64853
rect 130 64808 138 64842
rect 1572 64808 1580 64842
rect 130 64797 1580 64808
rect 130 64756 1580 64767
rect 130 64722 138 64756
rect 1572 64722 1580 64756
rect 130 64711 1580 64722
rect 130 64670 1580 64681
rect 130 64636 138 64670
rect 1572 64636 1580 64670
rect 130 64625 1580 64636
rect 130 64584 1580 64595
rect 130 64550 138 64584
rect 1572 64550 1580 64584
rect 130 64539 1580 64550
rect 130 64498 1580 64509
rect 130 64464 138 64498
rect 1572 64464 1580 64498
rect 130 64453 1580 64464
rect 130 64412 1580 64423
rect 130 64378 138 64412
rect 1572 64378 1580 64412
rect 130 64367 1580 64378
rect 130 64326 1580 64337
rect 130 64292 138 64326
rect 1572 64292 1580 64326
rect 130 64281 1580 64292
rect 130 64240 1580 64251
rect 130 64206 138 64240
rect 1572 64206 1580 64240
rect 130 64195 1580 64206
rect 130 64154 1580 64165
rect 130 64120 138 64154
rect 1572 64120 1580 64154
rect 130 64109 1580 64120
rect 130 64068 1580 64079
rect 130 64034 138 64068
rect 1572 64034 1580 64068
rect 130 64023 1580 64034
rect 130 63982 1580 63993
rect 130 63948 138 63982
rect 1572 63948 1580 63982
rect 130 63937 1580 63948
rect 130 63896 1580 63907
rect 130 63862 138 63896
rect 1572 63862 1580 63896
rect 130 63851 1580 63862
rect 130 63810 1580 63821
rect 130 63776 138 63810
rect 1572 63776 1580 63810
rect 130 63765 1580 63776
rect 130 63724 1580 63735
rect 130 63690 138 63724
rect 1572 63690 1580 63724
rect 130 63679 1580 63690
rect 130 63638 1580 63649
rect 130 63604 138 63638
rect 1572 63604 1580 63638
rect 130 63593 1580 63604
rect 130 63552 1580 63563
rect 130 63518 138 63552
rect 1572 63518 1580 63552
rect 130 63507 1580 63518
rect 130 63466 1580 63477
rect 130 63432 138 63466
rect 1572 63432 1580 63466
rect 130 63421 1580 63432
rect 130 63380 1580 63391
rect 130 63346 138 63380
rect 1572 63346 1580 63380
rect 130 63335 1580 63346
rect 130 63294 1580 63305
rect 130 63260 138 63294
rect 1572 63260 1580 63294
rect 130 63249 1580 63260
rect 130 63208 1580 63219
rect 130 63174 138 63208
rect 1572 63174 1580 63208
rect 130 63163 1580 63174
rect 130 63122 1580 63133
rect 130 63088 138 63122
rect 1572 63088 1580 63122
rect 130 63077 1580 63088
rect 130 63036 1580 63047
rect 130 63002 138 63036
rect 1572 63002 1580 63036
rect 130 62991 1580 63002
rect 130 62950 1580 62961
rect 130 62916 138 62950
rect 1572 62916 1580 62950
rect 130 62905 1580 62916
rect 130 62864 1580 62875
rect 130 62830 138 62864
rect 1572 62830 1580 62864
rect 130 62819 1580 62830
rect 130 62778 1580 62789
rect 130 62744 138 62778
rect 1572 62744 1580 62778
rect 130 62733 1580 62744
rect 130 62692 1580 62703
rect 130 62658 138 62692
rect 1572 62658 1580 62692
rect 130 62647 1580 62658
rect 130 62606 1580 62617
rect 130 62572 138 62606
rect 1572 62572 1580 62606
rect 130 62561 1580 62572
rect 130 62520 1580 62531
rect 130 62486 138 62520
rect 1572 62486 1580 62520
rect 130 62475 1580 62486
rect 130 62434 1580 62445
rect 130 62400 138 62434
rect 1572 62400 1580 62434
rect 130 62389 1580 62400
rect 130 62348 1580 62359
rect 130 62314 138 62348
rect 1572 62314 1580 62348
rect 130 62303 1580 62314
rect 130 62262 1580 62273
rect 130 62228 138 62262
rect 1572 62228 1580 62262
rect 130 62217 1580 62228
rect 130 62176 1580 62187
rect 130 62142 138 62176
rect 1572 62142 1580 62176
rect 130 62131 1580 62142
rect 130 62090 1580 62101
rect 130 62056 138 62090
rect 1572 62056 1580 62090
rect 130 62045 1580 62056
rect 130 62004 1580 62015
rect 130 61970 138 62004
rect 1572 61970 1580 62004
rect 130 61959 1580 61970
rect 130 61918 1580 61929
rect 130 61884 138 61918
rect 1572 61884 1580 61918
rect 130 61873 1580 61884
rect 130 61832 1580 61843
rect 130 61798 138 61832
rect 1572 61798 1580 61832
rect 130 61787 1580 61798
rect 130 61746 1580 61757
rect 130 61712 138 61746
rect 1572 61712 1580 61746
rect 130 61701 1580 61712
rect 130 61660 1580 61671
rect 130 61626 138 61660
rect 1572 61626 1580 61660
rect 130 61615 1580 61626
rect 130 61574 1580 61585
rect 130 61540 138 61574
rect 1572 61540 1580 61574
rect 130 61529 1580 61540
rect 130 61488 1580 61499
rect 130 61454 138 61488
rect 1572 61454 1580 61488
rect 130 61443 1580 61454
rect 130 61402 1580 61413
rect 130 61368 138 61402
rect 1572 61368 1580 61402
rect 130 61357 1580 61368
rect 130 61316 1580 61327
rect 130 61282 138 61316
rect 1572 61282 1580 61316
rect 130 61271 1580 61282
rect 130 61230 1580 61241
rect 130 61196 138 61230
rect 1572 61196 1580 61230
rect 130 61185 1580 61196
rect 130 61144 1580 61155
rect 130 61110 138 61144
rect 1572 61110 1580 61144
rect 130 61099 1580 61110
rect 130 61058 1580 61069
rect 130 61024 138 61058
rect 1572 61024 1580 61058
rect 130 61013 1580 61024
rect 130 60972 1580 60983
rect 130 60938 138 60972
rect 1572 60938 1580 60972
rect 130 60927 1580 60938
rect 130 60886 1580 60897
rect 130 60852 138 60886
rect 1572 60852 1580 60886
rect 130 60841 1580 60852
rect 130 60800 1580 60811
rect 130 60766 138 60800
rect 1572 60766 1580 60800
rect 130 60755 1580 60766
rect 130 60714 1580 60725
rect 130 60680 138 60714
rect 1572 60680 1580 60714
rect 130 60669 1580 60680
rect 130 60628 1580 60639
rect 130 60594 138 60628
rect 1572 60594 1580 60628
rect 130 60583 1580 60594
rect 130 60542 1580 60553
rect 130 60508 138 60542
rect 1572 60508 1580 60542
rect 130 60497 1580 60508
rect 130 60456 1580 60467
rect 130 60422 138 60456
rect 1572 60422 1580 60456
rect 130 60411 1580 60422
rect 130 60370 1580 60381
rect 130 60336 138 60370
rect 1572 60336 1580 60370
rect 130 60325 1580 60336
rect 130 60284 1580 60295
rect 130 60250 138 60284
rect 1572 60250 1580 60284
rect 130 60239 1580 60250
rect 130 60198 1580 60209
rect 130 60164 138 60198
rect 1572 60164 1580 60198
rect 130 60153 1580 60164
rect 130 60112 1580 60123
rect 130 60078 138 60112
rect 1572 60078 1580 60112
rect 130 60067 1580 60078
rect 130 60026 1580 60037
rect 130 59992 138 60026
rect 1572 59992 1580 60026
rect 130 59981 1580 59992
rect 130 59940 1580 59951
rect 130 59906 138 59940
rect 1572 59906 1580 59940
rect 130 59895 1580 59906
rect 130 59854 1580 59865
rect 130 59820 138 59854
rect 1572 59820 1580 59854
rect 130 59809 1580 59820
rect 130 59768 1580 59779
rect 130 59734 138 59768
rect 1572 59734 1580 59768
rect 130 59723 1580 59734
rect 130 59682 1580 59693
rect 130 59648 138 59682
rect 1572 59648 1580 59682
rect 130 59637 1580 59648
rect 130 59596 1580 59607
rect 130 59562 138 59596
rect 1572 59562 1580 59596
rect 130 59551 1580 59562
rect 130 59510 1580 59521
rect 130 59476 138 59510
rect 1572 59476 1580 59510
rect 130 59465 1580 59476
rect 130 59424 1580 59435
rect 130 59390 138 59424
rect 1572 59390 1580 59424
rect 130 59379 1580 59390
rect 130 59338 1580 59349
rect 130 59304 138 59338
rect 1572 59304 1580 59338
rect 130 59293 1580 59304
rect 130 59252 1580 59263
rect 130 59218 138 59252
rect 1572 59218 1580 59252
rect 130 59207 1580 59218
rect 130 59166 1580 59177
rect 130 59132 138 59166
rect 1572 59132 1580 59166
rect 130 59121 1580 59132
rect 130 59080 1580 59091
rect 130 59046 138 59080
rect 1572 59046 1580 59080
rect 130 59035 1580 59046
rect 130 58994 1580 59005
rect 130 58960 138 58994
rect 1572 58960 1580 58994
rect 130 58949 1580 58960
rect 130 58908 1580 58919
rect 130 58874 138 58908
rect 1572 58874 1580 58908
rect 130 58863 1580 58874
rect 130 58822 1580 58833
rect 130 58788 138 58822
rect 1572 58788 1580 58822
rect 130 58777 1580 58788
rect 130 58736 1580 58747
rect 130 58702 138 58736
rect 1572 58702 1580 58736
rect 130 58691 1580 58702
rect 130 58650 1580 58661
rect 130 58616 138 58650
rect 1572 58616 1580 58650
rect 130 58605 1580 58616
rect 130 58564 1580 58575
rect 130 58530 138 58564
rect 1572 58530 1580 58564
rect 130 58519 1580 58530
rect 130 58478 1580 58489
rect 130 58444 138 58478
rect 1572 58444 1580 58478
rect 130 58433 1580 58444
rect 130 58392 1580 58403
rect 130 58358 138 58392
rect 1572 58358 1580 58392
rect 130 58347 1580 58358
rect 130 58306 1580 58317
rect 130 58272 138 58306
rect 1572 58272 1580 58306
rect 130 58261 1580 58272
rect 130 58220 1580 58231
rect 130 58186 138 58220
rect 1572 58186 1580 58220
rect 130 58175 1580 58186
rect 130 58134 1580 58145
rect 130 58100 138 58134
rect 1572 58100 1580 58134
rect 130 58089 1580 58100
rect 130 58048 1580 58059
rect 130 58014 138 58048
rect 1572 58014 1580 58048
rect 130 58003 1580 58014
rect 130 57962 1580 57973
rect 130 57928 138 57962
rect 1572 57928 1580 57962
rect 130 57917 1580 57928
rect 130 57876 1580 57887
rect 130 57842 138 57876
rect 1572 57842 1580 57876
rect 130 57831 1580 57842
rect 130 57790 1580 57801
rect 130 57756 138 57790
rect 1572 57756 1580 57790
rect 130 57745 1580 57756
rect 130 57704 1580 57715
rect 130 57670 138 57704
rect 1572 57670 1580 57704
rect 130 57659 1580 57670
rect 130 57618 1580 57629
rect 130 57584 138 57618
rect 1572 57584 1580 57618
rect 130 57573 1580 57584
rect 130 57532 1580 57543
rect 130 57498 138 57532
rect 1572 57498 1580 57532
rect 130 57487 1580 57498
rect 130 57446 1580 57457
rect 130 57412 138 57446
rect 1572 57412 1580 57446
rect 130 57401 1580 57412
rect 130 57360 1580 57371
rect 130 57326 138 57360
rect 1572 57326 1580 57360
rect 130 57315 1580 57326
rect 130 57274 1580 57285
rect 130 57240 138 57274
rect 1572 57240 1580 57274
rect 130 57229 1580 57240
rect 130 57188 1580 57199
rect 130 57154 138 57188
rect 1572 57154 1580 57188
rect 130 57143 1580 57154
rect 130 57102 1580 57113
rect 130 57068 138 57102
rect 1572 57068 1580 57102
rect 130 57057 1580 57068
rect 130 57016 1580 57027
rect 130 56982 138 57016
rect 1572 56982 1580 57016
rect 130 56971 1580 56982
rect 130 56930 1580 56941
rect 130 56896 138 56930
rect 1572 56896 1580 56930
rect 130 56885 1580 56896
rect 130 56844 1580 56855
rect 130 56810 138 56844
rect 1572 56810 1580 56844
rect 130 56799 1580 56810
rect 130 56758 1580 56769
rect 130 56724 138 56758
rect 1572 56724 1580 56758
rect 130 56713 1580 56724
rect 130 56672 1580 56683
rect 130 56638 138 56672
rect 1572 56638 1580 56672
rect 130 56627 1580 56638
rect 130 56586 1580 56597
rect 130 56552 138 56586
rect 1572 56552 1580 56586
rect 130 56541 1580 56552
rect 130 56500 1580 56511
rect 130 56466 138 56500
rect 1572 56466 1580 56500
rect 130 56455 1580 56466
rect 130 56414 1580 56425
rect 130 56380 138 56414
rect 1572 56380 1580 56414
rect 130 56369 1580 56380
rect 130 56328 1580 56339
rect 130 56294 138 56328
rect 1572 56294 1580 56328
rect 130 56283 1580 56294
rect 130 56242 1580 56253
rect 130 56208 138 56242
rect 1572 56208 1580 56242
rect 130 56197 1580 56208
rect 130 56156 1580 56167
rect 130 56122 138 56156
rect 1572 56122 1580 56156
rect 130 56111 1580 56122
rect 130 56070 1580 56081
rect 130 56036 138 56070
rect 1572 56036 1580 56070
rect 130 56025 1580 56036
rect 130 55984 1580 55995
rect 130 55950 138 55984
rect 1572 55950 1580 55984
rect 130 55939 1580 55950
rect 130 55898 1580 55909
rect 130 55864 138 55898
rect 1572 55864 1580 55898
rect 130 55853 1580 55864
rect 130 55812 1580 55823
rect 130 55778 138 55812
rect 1572 55778 1580 55812
rect 130 55767 1580 55778
rect 130 55726 1580 55737
rect 130 55692 138 55726
rect 1572 55692 1580 55726
rect 130 55681 1580 55692
rect 130 55640 1580 55651
rect 130 55606 138 55640
rect 1572 55606 1580 55640
rect 130 55595 1580 55606
rect 130 55554 1580 55565
rect 130 55520 138 55554
rect 1572 55520 1580 55554
rect 130 55509 1580 55520
rect 130 55468 1580 55479
rect 130 55434 138 55468
rect 1572 55434 1580 55468
rect 130 55423 1580 55434
rect 130 55382 1580 55393
rect 130 55348 138 55382
rect 1572 55348 1580 55382
rect 130 55337 1580 55348
rect 130 55296 1580 55307
rect 130 55262 138 55296
rect 1572 55262 1580 55296
rect 130 55251 1580 55262
rect 130 55210 1580 55221
rect 130 55176 138 55210
rect 1572 55176 1580 55210
rect 130 55165 1580 55176
rect 130 55124 1580 55135
rect 130 55090 138 55124
rect 1572 55090 1580 55124
rect 130 55079 1580 55090
rect 130 55038 1580 55049
rect 130 55004 138 55038
rect 1572 55004 1580 55038
rect 130 54993 1580 55004
rect 130 54952 1580 54963
rect 130 54918 138 54952
rect 1572 54918 1580 54952
rect 130 54907 1580 54918
rect 130 54866 1580 54877
rect 130 54832 138 54866
rect 1572 54832 1580 54866
rect 130 54821 1580 54832
rect 130 54780 1580 54791
rect 130 54746 138 54780
rect 1572 54746 1580 54780
rect 130 54735 1580 54746
rect 130 54694 1580 54705
rect 130 54660 138 54694
rect 1572 54660 1580 54694
rect 130 54649 1580 54660
rect 130 54608 1580 54619
rect 130 54574 138 54608
rect 1572 54574 1580 54608
rect 130 54563 1580 54574
rect 130 54522 1580 54533
rect 130 54488 138 54522
rect 1572 54488 1580 54522
rect 130 54477 1580 54488
rect 130 54436 1580 54447
rect 130 54402 138 54436
rect 1572 54402 1580 54436
rect 130 54391 1580 54402
rect 130 54350 1580 54361
rect 130 54316 138 54350
rect 1572 54316 1580 54350
rect 130 54305 1580 54316
rect 130 54264 1580 54275
rect 130 54230 138 54264
rect 1572 54230 1580 54264
rect 130 54219 1580 54230
rect 130 54178 1580 54189
rect 130 54144 138 54178
rect 1572 54144 1580 54178
rect 130 54133 1580 54144
rect 130 54092 1580 54103
rect 130 54058 138 54092
rect 1572 54058 1580 54092
rect 130 54047 1580 54058
rect 130 54006 1580 54017
rect 130 53972 138 54006
rect 1572 53972 1580 54006
rect 130 53961 1580 53972
rect 130 53920 1580 53931
rect 130 53886 138 53920
rect 1572 53886 1580 53920
rect 130 53875 1580 53886
rect 130 53834 1580 53845
rect 130 53800 138 53834
rect 1572 53800 1580 53834
rect 130 53789 1580 53800
rect 130 53748 1580 53759
rect 130 53714 138 53748
rect 1572 53714 1580 53748
rect 130 53703 1580 53714
rect 130 53662 1580 53673
rect 130 53628 138 53662
rect 1572 53628 1580 53662
rect 130 53617 1580 53628
rect 130 53576 1580 53587
rect 130 53542 138 53576
rect 1572 53542 1580 53576
rect 130 53531 1580 53542
rect 130 53490 1580 53501
rect 130 53456 138 53490
rect 1572 53456 1580 53490
rect 130 53445 1580 53456
rect 130 53404 1580 53415
rect 130 53370 138 53404
rect 1572 53370 1580 53404
rect 130 53359 1580 53370
rect 130 53318 1580 53329
rect 130 53284 138 53318
rect 1572 53284 1580 53318
rect 130 53273 1580 53284
rect 130 53232 1580 53243
rect 130 53198 138 53232
rect 1572 53198 1580 53232
rect 130 53187 1580 53198
rect 130 53146 1580 53157
rect 130 53112 138 53146
rect 1572 53112 1580 53146
rect 130 53101 1580 53112
rect 130 53060 1580 53071
rect 130 53026 138 53060
rect 1572 53026 1580 53060
rect 130 53015 1580 53026
rect 130 52974 1580 52985
rect 130 52940 138 52974
rect 1572 52940 1580 52974
rect 130 52929 1580 52940
rect 130 52888 1580 52899
rect 130 52854 138 52888
rect 1572 52854 1580 52888
rect 130 52843 1580 52854
rect 130 52802 1580 52813
rect 130 52768 138 52802
rect 1572 52768 1580 52802
rect 130 52757 1580 52768
rect 130 52716 1580 52727
rect 130 52682 138 52716
rect 1572 52682 1580 52716
rect 130 52671 1580 52682
rect 130 52630 1580 52641
rect 130 52596 138 52630
rect 1572 52596 1580 52630
rect 130 52585 1580 52596
rect 130 52544 1580 52555
rect 130 52510 138 52544
rect 1572 52510 1580 52544
rect 130 52499 1580 52510
rect 130 52458 1580 52469
rect 130 52424 138 52458
rect 1572 52424 1580 52458
rect 130 52413 1580 52424
rect 130 52372 1580 52383
rect 130 52338 138 52372
rect 1572 52338 1580 52372
rect 130 52327 1580 52338
rect 130 52286 1580 52297
rect 130 52252 138 52286
rect 1572 52252 1580 52286
rect 130 52241 1580 52252
rect 130 52200 1580 52211
rect 130 52166 138 52200
rect 1572 52166 1580 52200
rect 130 52155 1580 52166
rect 130 52114 1580 52125
rect 130 52080 138 52114
rect 1572 52080 1580 52114
rect 130 52069 1580 52080
rect 130 52028 1580 52039
rect 130 51994 138 52028
rect 1572 51994 1580 52028
rect 130 51983 1580 51994
rect 130 51942 1580 51953
rect 130 51908 138 51942
rect 1572 51908 1580 51942
rect 130 51897 1580 51908
rect 130 51856 1580 51867
rect 130 51822 138 51856
rect 1572 51822 1580 51856
rect 130 51811 1580 51822
rect 130 51770 1580 51781
rect 130 51736 138 51770
rect 1572 51736 1580 51770
rect 130 51725 1580 51736
rect 130 51684 1580 51695
rect 130 51650 138 51684
rect 1572 51650 1580 51684
rect 130 51639 1580 51650
rect 130 51598 1580 51609
rect 130 51564 138 51598
rect 1572 51564 1580 51598
rect 130 51553 1580 51564
rect 130 51512 1580 51523
rect 130 51478 138 51512
rect 1572 51478 1580 51512
rect 130 51467 1580 51478
rect 130 51426 1580 51437
rect 130 51392 138 51426
rect 1572 51392 1580 51426
rect 130 51381 1580 51392
rect 130 51340 1580 51351
rect 130 51306 138 51340
rect 1572 51306 1580 51340
rect 130 51295 1580 51306
rect 130 51254 1580 51265
rect 130 51220 138 51254
rect 1572 51220 1580 51254
rect 130 51209 1580 51220
rect 130 51168 1580 51179
rect 130 51134 138 51168
rect 1572 51134 1580 51168
rect 130 51123 1580 51134
rect 130 51082 1580 51093
rect 130 51048 138 51082
rect 1572 51048 1580 51082
rect 130 51037 1580 51048
rect 130 50996 1580 51007
rect 130 50962 138 50996
rect 1572 50962 1580 50996
rect 130 50951 1580 50962
rect 130 50910 1580 50921
rect 130 50876 138 50910
rect 1572 50876 1580 50910
rect 130 50865 1580 50876
rect 130 50824 1580 50835
rect 130 50790 138 50824
rect 1572 50790 1580 50824
rect 130 50779 1580 50790
rect 130 50738 1580 50749
rect 130 50704 138 50738
rect 1572 50704 1580 50738
rect 130 50693 1580 50704
rect 130 50652 1580 50663
rect 130 50618 138 50652
rect 1572 50618 1580 50652
rect 130 50607 1580 50618
rect 130 50566 1580 50577
rect 130 50532 138 50566
rect 1572 50532 1580 50566
rect 130 50521 1580 50532
rect 130 50480 1580 50491
rect 130 50446 138 50480
rect 1572 50446 1580 50480
rect 130 50435 1580 50446
rect 130 50394 1580 50405
rect 130 50360 138 50394
rect 1572 50360 1580 50394
rect 130 50349 1580 50360
rect 130 50308 1580 50319
rect 130 50274 138 50308
rect 1572 50274 1580 50308
rect 130 50263 1580 50274
rect 130 50222 1580 50233
rect 130 50188 138 50222
rect 1572 50188 1580 50222
rect 130 50177 1580 50188
rect 130 50136 1580 50147
rect 130 50102 138 50136
rect 1572 50102 1580 50136
rect 130 50091 1580 50102
rect 130 50050 1580 50061
rect 130 50016 138 50050
rect 1572 50016 1580 50050
rect 130 50005 1580 50016
rect 130 49964 1580 49975
rect 130 49930 138 49964
rect 1572 49930 1580 49964
rect 130 49919 1580 49930
rect 130 49878 1580 49889
rect 130 49844 138 49878
rect 1572 49844 1580 49878
rect 130 49833 1580 49844
rect 130 49792 1580 49803
rect 130 49758 138 49792
rect 1572 49758 1580 49792
rect 130 49747 1580 49758
rect 130 49706 1580 49717
rect 130 49672 138 49706
rect 1572 49672 1580 49706
rect 130 49661 1580 49672
rect 130 49620 1580 49631
rect 130 49586 138 49620
rect 1572 49586 1580 49620
rect 130 49575 1580 49586
rect 130 49534 1580 49545
rect 130 49500 138 49534
rect 1572 49500 1580 49534
rect 130 49489 1580 49500
rect 130 49448 1580 49459
rect 130 49414 138 49448
rect 1572 49414 1580 49448
rect 130 49403 1580 49414
rect 130 49362 1580 49373
rect 130 49328 138 49362
rect 1572 49328 1580 49362
rect 130 49317 1580 49328
rect 130 49276 1580 49287
rect 130 49242 138 49276
rect 1572 49242 1580 49276
rect 130 49231 1580 49242
rect 130 49190 1580 49201
rect 130 49156 138 49190
rect 1572 49156 1580 49190
rect 130 49145 1580 49156
rect 130 49104 1580 49115
rect 130 49070 138 49104
rect 1572 49070 1580 49104
rect 130 49059 1580 49070
rect 130 49018 1580 49029
rect 130 48984 138 49018
rect 1572 48984 1580 49018
rect 130 48973 1580 48984
rect 130 48932 1580 48943
rect 130 48898 138 48932
rect 1572 48898 1580 48932
rect 130 48887 1580 48898
rect 130 48846 1580 48857
rect 130 48812 138 48846
rect 1572 48812 1580 48846
rect 130 48801 1580 48812
rect 130 48760 1580 48771
rect 130 48726 138 48760
rect 1572 48726 1580 48760
rect 130 48715 1580 48726
rect 130 48674 1580 48685
rect 130 48640 138 48674
rect 1572 48640 1580 48674
rect 130 48629 1580 48640
rect 130 48588 1580 48599
rect 130 48554 138 48588
rect 1572 48554 1580 48588
rect 130 48543 1580 48554
rect 130 48502 1580 48513
rect 130 48468 138 48502
rect 1572 48468 1580 48502
rect 130 48457 1580 48468
rect 130 48416 1580 48427
rect 130 48382 138 48416
rect 1572 48382 1580 48416
rect 130 48371 1580 48382
rect 130 48330 1580 48341
rect 130 48296 138 48330
rect 1572 48296 1580 48330
rect 130 48285 1580 48296
rect 130 48244 1580 48255
rect 130 48210 138 48244
rect 1572 48210 1580 48244
rect 130 48199 1580 48210
rect 130 48158 1580 48169
rect 130 48124 138 48158
rect 1572 48124 1580 48158
rect 130 48113 1580 48124
rect 130 48072 1580 48083
rect 130 48038 138 48072
rect 1572 48038 1580 48072
rect 130 48027 1580 48038
rect 130 47986 1580 47997
rect 130 47952 138 47986
rect 1572 47952 1580 47986
rect 130 47941 1580 47952
rect 130 47900 1580 47911
rect 130 47866 138 47900
rect 1572 47866 1580 47900
rect 130 47855 1580 47866
rect 130 47814 1580 47825
rect 130 47780 138 47814
rect 1572 47780 1580 47814
rect 130 47769 1580 47780
rect 130 47728 1580 47739
rect 130 47694 138 47728
rect 1572 47694 1580 47728
rect 130 47683 1580 47694
rect 130 47642 1580 47653
rect 130 47608 138 47642
rect 1572 47608 1580 47642
rect 130 47597 1580 47608
rect 130 47556 1580 47567
rect 130 47522 138 47556
rect 1572 47522 1580 47556
rect 130 47511 1580 47522
rect 130 47470 1580 47481
rect 130 47436 138 47470
rect 1572 47436 1580 47470
rect 130 47425 1580 47436
rect 130 47384 1580 47395
rect 130 47350 138 47384
rect 1572 47350 1580 47384
rect 130 47339 1580 47350
rect 130 47298 1580 47309
rect 130 47264 138 47298
rect 1572 47264 1580 47298
rect 130 47253 1580 47264
rect 130 47212 1580 47223
rect 130 47178 138 47212
rect 1572 47178 1580 47212
rect 130 47167 1580 47178
rect 130 47126 1580 47137
rect 130 47092 138 47126
rect 1572 47092 1580 47126
rect 130 47081 1580 47092
rect 130 47040 1580 47051
rect 130 47006 138 47040
rect 1572 47006 1580 47040
rect 130 46995 1580 47006
rect 130 46954 1580 46965
rect 130 46920 138 46954
rect 1572 46920 1580 46954
rect 130 46909 1580 46920
rect 130 46868 1580 46879
rect 130 46834 138 46868
rect 1572 46834 1580 46868
rect 130 46823 1580 46834
rect 130 46782 1580 46793
rect 130 46748 138 46782
rect 1572 46748 1580 46782
rect 130 46737 1580 46748
rect 130 46696 1580 46707
rect 130 46662 138 46696
rect 1572 46662 1580 46696
rect 130 46651 1580 46662
rect 130 46610 1580 46621
rect 130 46576 138 46610
rect 1572 46576 1580 46610
rect 130 46565 1580 46576
rect 130 46524 1580 46535
rect 130 46490 138 46524
rect 1572 46490 1580 46524
rect 130 46479 1580 46490
rect 130 46438 1580 46449
rect 130 46404 138 46438
rect 1572 46404 1580 46438
rect 130 46393 1580 46404
rect 130 46352 1580 46363
rect 130 46318 138 46352
rect 1572 46318 1580 46352
rect 130 46307 1580 46318
rect 130 46266 1580 46277
rect 130 46232 138 46266
rect 1572 46232 1580 46266
rect 130 46221 1580 46232
rect 130 46180 1580 46191
rect 130 46146 138 46180
rect 1572 46146 1580 46180
rect 130 46135 1580 46146
rect 130 46094 1580 46105
rect 130 46060 138 46094
rect 1572 46060 1580 46094
rect 130 46049 1580 46060
rect 130 46008 1580 46019
rect 130 45974 138 46008
rect 1572 45974 1580 46008
rect 130 45963 1580 45974
rect 130 45922 1580 45933
rect 130 45888 138 45922
rect 1572 45888 1580 45922
rect 130 45877 1580 45888
rect 130 45836 1580 45847
rect 130 45802 138 45836
rect 1572 45802 1580 45836
rect 130 45791 1580 45802
rect 130 45750 1580 45761
rect 130 45716 138 45750
rect 1572 45716 1580 45750
rect 130 45705 1580 45716
rect 130 45664 1580 45675
rect 130 45630 138 45664
rect 1572 45630 1580 45664
rect 130 45619 1580 45630
rect 130 45578 1580 45589
rect 130 45544 138 45578
rect 1572 45544 1580 45578
rect 130 45533 1580 45544
rect 130 45492 1580 45503
rect 130 45458 138 45492
rect 1572 45458 1580 45492
rect 130 45447 1580 45458
rect 130 45406 1580 45417
rect 130 45372 138 45406
rect 1572 45372 1580 45406
rect 130 45361 1580 45372
rect 130 45320 1580 45331
rect 130 45286 138 45320
rect 1572 45286 1580 45320
rect 130 45275 1580 45286
rect 130 45234 1580 45245
rect 130 45200 138 45234
rect 1572 45200 1580 45234
rect 130 45189 1580 45200
rect 130 45148 1580 45159
rect 130 45114 138 45148
rect 1572 45114 1580 45148
rect 130 45103 1580 45114
rect 130 45062 1580 45073
rect 130 45028 138 45062
rect 1572 45028 1580 45062
rect 130 45017 1580 45028
rect 130 44976 1580 44987
rect 130 44942 138 44976
rect 1572 44942 1580 44976
rect 130 44931 1580 44942
rect 130 44890 1580 44901
rect 130 44856 138 44890
rect 1572 44856 1580 44890
rect 130 44845 1580 44856
rect 130 44804 1580 44815
rect 130 44770 138 44804
rect 1572 44770 1580 44804
rect 130 44759 1580 44770
rect 130 44718 1580 44729
rect 130 44684 138 44718
rect 1572 44684 1580 44718
rect 130 44673 1580 44684
rect 130 44632 1580 44643
rect 130 44598 138 44632
rect 1572 44598 1580 44632
rect 130 44587 1580 44598
rect 130 44546 1580 44557
rect 130 44512 138 44546
rect 1572 44512 1580 44546
rect 130 44501 1580 44512
rect 130 44460 1580 44471
rect 130 44426 138 44460
rect 1572 44426 1580 44460
rect 130 44415 1580 44426
rect 130 44374 1580 44385
rect 130 44340 138 44374
rect 1572 44340 1580 44374
rect 130 44329 1580 44340
rect 130 44288 1580 44299
rect 130 44254 138 44288
rect 1572 44254 1580 44288
rect 130 44243 1580 44254
rect 130 44202 1580 44213
rect 130 44168 138 44202
rect 1572 44168 1580 44202
rect 130 44157 1580 44168
rect 130 44116 1580 44127
rect 130 44082 138 44116
rect 1572 44082 1580 44116
rect 130 44071 1580 44082
rect 130 44030 1580 44041
rect 130 43996 138 44030
rect 1572 43996 1580 44030
rect 130 43985 1580 43996
rect 130 43944 1580 43955
rect 130 43910 138 43944
rect 1572 43910 1580 43944
rect 130 43899 1580 43910
rect 130 43858 1580 43869
rect 130 43824 138 43858
rect 1572 43824 1580 43858
rect 130 43813 1580 43824
rect 130 43772 1580 43783
rect 130 43738 138 43772
rect 1572 43738 1580 43772
rect 130 43727 1580 43738
rect 130 43686 1580 43697
rect 130 43652 138 43686
rect 1572 43652 1580 43686
rect 130 43641 1580 43652
rect 130 43600 1580 43611
rect 130 43566 138 43600
rect 1572 43566 1580 43600
rect 130 43555 1580 43566
rect 130 43514 1580 43525
rect 130 43480 138 43514
rect 1572 43480 1580 43514
rect 130 43469 1580 43480
rect 130 43428 1580 43439
rect 130 43394 138 43428
rect 1572 43394 1580 43428
rect 130 43383 1580 43394
rect 130 43342 1580 43353
rect 130 43308 138 43342
rect 1572 43308 1580 43342
rect 130 43297 1580 43308
rect 130 43256 1580 43267
rect 130 43222 138 43256
rect 1572 43222 1580 43256
rect 130 43211 1580 43222
rect 130 43170 1580 43181
rect 130 43136 138 43170
rect 1572 43136 1580 43170
rect 130 43125 1580 43136
rect 130 43084 1580 43095
rect 130 43050 138 43084
rect 1572 43050 1580 43084
rect 130 43039 1580 43050
rect 130 42998 1580 43009
rect 130 42964 138 42998
rect 1572 42964 1580 42998
rect 130 42953 1580 42964
rect 130 42912 1580 42923
rect 130 42878 138 42912
rect 1572 42878 1580 42912
rect 130 42867 1580 42878
rect 130 42826 1580 42837
rect 130 42792 138 42826
rect 1572 42792 1580 42826
rect 130 42781 1580 42792
rect 130 42740 1580 42751
rect 130 42706 138 42740
rect 1572 42706 1580 42740
rect 130 42695 1580 42706
rect 130 42654 1580 42665
rect 130 42620 138 42654
rect 1572 42620 1580 42654
rect 130 42609 1580 42620
rect 130 42568 1580 42579
rect 130 42534 138 42568
rect 1572 42534 1580 42568
rect 130 42523 1580 42534
rect 130 42482 1580 42493
rect 130 42448 138 42482
rect 1572 42448 1580 42482
rect 130 42437 1580 42448
rect 130 42396 1580 42407
rect 130 42362 138 42396
rect 1572 42362 1580 42396
rect 130 42351 1580 42362
rect 130 42310 1580 42321
rect 130 42276 138 42310
rect 1572 42276 1580 42310
rect 130 42265 1580 42276
rect 130 42224 1580 42235
rect 130 42190 138 42224
rect 1572 42190 1580 42224
rect 130 42179 1580 42190
rect 130 42138 1580 42149
rect 130 42104 138 42138
rect 1572 42104 1580 42138
rect 130 42093 1580 42104
rect 130 42052 1580 42063
rect 130 42018 138 42052
rect 1572 42018 1580 42052
rect 130 42007 1580 42018
rect 130 41966 1580 41977
rect 130 41932 138 41966
rect 1572 41932 1580 41966
rect 130 41921 1580 41932
rect 130 41880 1580 41891
rect 130 41846 138 41880
rect 1572 41846 1580 41880
rect 130 41835 1580 41846
rect 130 41794 1580 41805
rect 130 41760 138 41794
rect 1572 41760 1580 41794
rect 130 41749 1580 41760
rect 130 41708 1580 41719
rect 130 41674 138 41708
rect 1572 41674 1580 41708
rect 130 41663 1580 41674
rect 130 41622 1580 41633
rect 130 41588 138 41622
rect 1572 41588 1580 41622
rect 130 41577 1580 41588
rect 130 41536 1580 41547
rect 130 41502 138 41536
rect 1572 41502 1580 41536
rect 130 41491 1580 41502
rect 130 41450 1580 41461
rect 130 41416 138 41450
rect 1572 41416 1580 41450
rect 130 41405 1580 41416
rect 130 41364 1580 41375
rect 130 41330 138 41364
rect 1572 41330 1580 41364
rect 130 41319 1580 41330
rect 130 41278 1580 41289
rect 130 41244 138 41278
rect 1572 41244 1580 41278
rect 130 41233 1580 41244
rect 130 41192 1580 41203
rect 130 41158 138 41192
rect 1572 41158 1580 41192
rect 130 41147 1580 41158
rect 130 41106 1580 41117
rect 130 41072 138 41106
rect 1572 41072 1580 41106
rect 130 41061 1580 41072
rect 130 41020 1580 41031
rect 130 40986 138 41020
rect 1572 40986 1580 41020
rect 130 40975 1580 40986
rect 130 40934 1580 40945
rect 130 40900 138 40934
rect 1572 40900 1580 40934
rect 130 40889 1580 40900
rect 130 40848 1580 40859
rect 130 40814 138 40848
rect 1572 40814 1580 40848
rect 130 40803 1580 40814
rect 130 40762 1580 40773
rect 130 40728 138 40762
rect 1572 40728 1580 40762
rect 130 40717 1580 40728
rect 130 40676 1580 40687
rect 130 40642 138 40676
rect 1572 40642 1580 40676
rect 130 40631 1580 40642
rect 130 40590 1580 40601
rect 130 40556 138 40590
rect 1572 40556 1580 40590
rect 130 40545 1580 40556
rect 130 40504 1580 40515
rect 130 40470 138 40504
rect 1572 40470 1580 40504
rect 130 40459 1580 40470
rect 130 40418 1580 40429
rect 130 40384 138 40418
rect 1572 40384 1580 40418
rect 130 40373 1580 40384
rect 130 40332 1580 40343
rect 130 40298 138 40332
rect 1572 40298 1580 40332
rect 130 40287 1580 40298
rect 130 40246 1580 40257
rect 130 40212 138 40246
rect 1572 40212 1580 40246
rect 130 40201 1580 40212
rect 130 40160 1580 40171
rect 130 40126 138 40160
rect 1572 40126 1580 40160
rect 130 40115 1580 40126
rect 130 40074 1580 40085
rect 130 40040 138 40074
rect 1572 40040 1580 40074
rect 130 40029 1580 40040
rect 130 39988 1580 39999
rect 130 39954 138 39988
rect 1572 39954 1580 39988
rect 130 39943 1580 39954
rect 130 39902 1580 39913
rect 130 39868 138 39902
rect 1572 39868 1580 39902
rect 130 39857 1580 39868
rect 130 39816 1580 39827
rect 130 39782 138 39816
rect 1572 39782 1580 39816
rect 130 39771 1580 39782
rect 130 39730 1580 39741
rect 130 39696 138 39730
rect 1572 39696 1580 39730
rect 130 39685 1580 39696
rect 130 39644 1580 39655
rect 130 39610 138 39644
rect 1572 39610 1580 39644
rect 130 39599 1580 39610
rect 130 39558 1580 39569
rect 130 39524 138 39558
rect 1572 39524 1580 39558
rect 130 39513 1580 39524
rect 130 39472 1580 39483
rect 130 39438 138 39472
rect 1572 39438 1580 39472
rect 130 39427 1580 39438
rect 130 39386 1580 39397
rect 130 39352 138 39386
rect 1572 39352 1580 39386
rect 130 39341 1580 39352
rect 130 39300 1580 39311
rect 130 39266 138 39300
rect 1572 39266 1580 39300
rect 130 39255 1580 39266
rect 130 39214 1580 39225
rect 130 39180 138 39214
rect 1572 39180 1580 39214
rect 130 39169 1580 39180
rect 130 39128 1580 39139
rect 130 39094 138 39128
rect 1572 39094 1580 39128
rect 130 39083 1580 39094
rect 130 39042 1580 39053
rect 130 39008 138 39042
rect 1572 39008 1580 39042
rect 130 38997 1580 39008
rect 130 38956 1580 38967
rect 130 38922 138 38956
rect 1572 38922 1580 38956
rect 130 38911 1580 38922
rect 130 38870 1580 38881
rect 130 38836 138 38870
rect 1572 38836 1580 38870
rect 130 38825 1580 38836
rect 130 38784 1580 38795
rect 130 38750 138 38784
rect 1572 38750 1580 38784
rect 130 38739 1580 38750
rect 130 38698 1580 38709
rect 130 38664 138 38698
rect 1572 38664 1580 38698
rect 130 38653 1580 38664
rect 130 38612 1580 38623
rect 130 38578 138 38612
rect 1572 38578 1580 38612
rect 130 38567 1580 38578
rect 130 38526 1580 38537
rect 130 38492 138 38526
rect 1572 38492 1580 38526
rect 130 38481 1580 38492
rect 130 38440 1580 38451
rect 130 38406 138 38440
rect 1572 38406 1580 38440
rect 130 38395 1580 38406
rect 130 38354 1580 38365
rect 130 38320 138 38354
rect 1572 38320 1580 38354
rect 130 38309 1580 38320
rect 130 38268 1580 38279
rect 130 38234 138 38268
rect 1572 38234 1580 38268
rect 130 38223 1580 38234
rect 130 38182 1580 38193
rect 130 38148 138 38182
rect 1572 38148 1580 38182
rect 130 38137 1580 38148
rect 130 38096 1580 38107
rect 130 38062 138 38096
rect 1572 38062 1580 38096
rect 130 38051 1580 38062
rect 130 38010 1580 38021
rect 130 37976 138 38010
rect 1572 37976 1580 38010
rect 130 37965 1580 37976
rect 130 37924 1580 37935
rect 130 37890 138 37924
rect 1572 37890 1580 37924
rect 130 37879 1580 37890
rect 130 37838 1580 37849
rect 130 37804 138 37838
rect 1572 37804 1580 37838
rect 130 37793 1580 37804
rect 130 37752 1580 37763
rect 130 37718 138 37752
rect 1572 37718 1580 37752
rect 130 37707 1580 37718
rect 130 37666 1580 37677
rect 130 37632 138 37666
rect 1572 37632 1580 37666
rect 130 37621 1580 37632
rect 130 37580 1580 37591
rect 130 37546 138 37580
rect 1572 37546 1580 37580
rect 130 37535 1580 37546
rect 130 37494 1580 37505
rect 130 37460 138 37494
rect 1572 37460 1580 37494
rect 130 37449 1580 37460
rect 130 37408 1580 37419
rect 130 37374 138 37408
rect 1572 37374 1580 37408
rect 130 37363 1580 37374
rect 130 37322 1580 37333
rect 130 37288 138 37322
rect 1572 37288 1580 37322
rect 130 37277 1580 37288
rect 130 37236 1580 37247
rect 130 37202 138 37236
rect 1572 37202 1580 37236
rect 130 37191 1580 37202
rect 130 37150 1580 37161
rect 130 37116 138 37150
rect 1572 37116 1580 37150
rect 130 37105 1580 37116
rect 130 37064 1580 37075
rect 130 37030 138 37064
rect 1572 37030 1580 37064
rect 130 37019 1580 37030
rect 130 36978 1580 36989
rect 130 36944 138 36978
rect 1572 36944 1580 36978
rect 130 36933 1580 36944
rect 130 36892 1580 36903
rect 130 36858 138 36892
rect 1572 36858 1580 36892
rect 130 36847 1580 36858
rect 130 36806 1580 36817
rect 130 36772 138 36806
rect 1572 36772 1580 36806
rect 130 36761 1580 36772
rect 130 36720 1580 36731
rect 130 36686 138 36720
rect 1572 36686 1580 36720
rect 130 36675 1580 36686
rect 130 36634 1580 36645
rect 130 36600 138 36634
rect 1572 36600 1580 36634
rect 130 36589 1580 36600
rect 130 36548 1580 36559
rect 130 36514 138 36548
rect 1572 36514 1580 36548
rect 130 36503 1580 36514
rect 130 36462 1580 36473
rect 130 36428 138 36462
rect 1572 36428 1580 36462
rect 130 36417 1580 36428
rect 130 36376 1580 36387
rect 130 36342 138 36376
rect 1572 36342 1580 36376
rect 130 36331 1580 36342
rect 130 36290 1580 36301
rect 130 36256 138 36290
rect 1572 36256 1580 36290
rect 130 36245 1580 36256
rect 130 36204 1580 36215
rect 130 36170 138 36204
rect 1572 36170 1580 36204
rect 130 36159 1580 36170
rect 130 36118 1580 36129
rect 130 36084 138 36118
rect 1572 36084 1580 36118
rect 130 36073 1580 36084
rect 130 36032 1580 36043
rect 130 35998 138 36032
rect 1572 35998 1580 36032
rect 130 35987 1580 35998
rect 130 35946 1580 35957
rect 130 35912 138 35946
rect 1572 35912 1580 35946
rect 130 35901 1580 35912
rect 130 35860 1580 35871
rect 130 35826 138 35860
rect 1572 35826 1580 35860
rect 130 35815 1580 35826
rect 130 35774 1580 35785
rect 130 35740 138 35774
rect 1572 35740 1580 35774
rect 130 35729 1580 35740
rect 130 35688 1580 35699
rect 130 35654 138 35688
rect 1572 35654 1580 35688
rect 130 35643 1580 35654
rect 130 35602 1580 35613
rect 130 35568 138 35602
rect 1572 35568 1580 35602
rect 130 35557 1580 35568
rect 130 35516 1580 35527
rect 130 35482 138 35516
rect 1572 35482 1580 35516
rect 130 35471 1580 35482
rect 130 35430 1580 35441
rect 130 35396 138 35430
rect 1572 35396 1580 35430
rect 130 35385 1580 35396
rect 130 35344 1580 35355
rect 130 35310 138 35344
rect 1572 35310 1580 35344
rect 130 35299 1580 35310
rect 130 35258 1580 35269
rect 130 35224 138 35258
rect 1572 35224 1580 35258
rect 130 35213 1580 35224
rect 130 35172 1580 35183
rect 130 35138 138 35172
rect 1572 35138 1580 35172
rect 130 35127 1580 35138
rect 130 35086 1580 35097
rect 130 35052 138 35086
rect 1572 35052 1580 35086
rect 130 35041 1580 35052
rect 130 35000 1580 35011
rect 130 34966 138 35000
rect 1572 34966 1580 35000
rect 130 34955 1580 34966
rect 130 34914 1580 34925
rect 130 34880 138 34914
rect 1572 34880 1580 34914
rect 130 34869 1580 34880
rect 130 34828 1580 34839
rect 130 34794 138 34828
rect 1572 34794 1580 34828
rect 130 34783 1580 34794
rect 130 34742 1580 34753
rect 130 34708 138 34742
rect 1572 34708 1580 34742
rect 130 34697 1580 34708
rect 130 34656 1580 34667
rect 130 34622 138 34656
rect 1572 34622 1580 34656
rect 130 34611 1580 34622
rect 130 34570 1580 34581
rect 130 34536 138 34570
rect 1572 34536 1580 34570
rect 130 34525 1580 34536
rect 130 34484 1580 34495
rect 130 34450 138 34484
rect 1572 34450 1580 34484
rect 130 34439 1580 34450
rect 130 34398 1580 34409
rect 130 34364 138 34398
rect 1572 34364 1580 34398
rect 130 34353 1580 34364
rect 130 34312 1580 34323
rect 130 34278 138 34312
rect 1572 34278 1580 34312
rect 130 34267 1580 34278
rect 130 34226 1580 34237
rect 130 34192 138 34226
rect 1572 34192 1580 34226
rect 130 34181 1580 34192
rect 130 34140 1580 34151
rect 130 34106 138 34140
rect 1572 34106 1580 34140
rect 130 34095 1580 34106
rect 130 34054 1580 34065
rect 130 34020 138 34054
rect 1572 34020 1580 34054
rect 130 34009 1580 34020
rect 130 33968 1580 33979
rect 130 33934 138 33968
rect 1572 33934 1580 33968
rect 130 33923 1580 33934
rect 130 33882 1580 33893
rect 130 33848 138 33882
rect 1572 33848 1580 33882
rect 130 33837 1580 33848
rect 130 33796 1580 33807
rect 130 33762 138 33796
rect 1572 33762 1580 33796
rect 130 33751 1580 33762
rect 130 33710 1580 33721
rect 130 33676 138 33710
rect 1572 33676 1580 33710
rect 130 33665 1580 33676
rect 130 33624 1580 33635
rect 130 33590 138 33624
rect 1572 33590 1580 33624
rect 130 33579 1580 33590
rect 130 33538 1580 33549
rect 130 33504 138 33538
rect 1572 33504 1580 33538
rect 130 33493 1580 33504
rect 130 33452 1580 33463
rect 130 33418 138 33452
rect 1572 33418 1580 33452
rect 130 33407 1580 33418
rect 130 33366 1580 33377
rect 130 33332 138 33366
rect 1572 33332 1580 33366
rect 130 33321 1580 33332
rect 130 33280 1580 33291
rect 130 33246 138 33280
rect 1572 33246 1580 33280
rect 130 33235 1580 33246
rect 130 33194 1580 33205
rect 130 33160 138 33194
rect 1572 33160 1580 33194
rect 130 33149 1580 33160
rect 130 33108 1580 33119
rect 130 33074 138 33108
rect 1572 33074 1580 33108
rect 130 33063 1580 33074
rect 130 33022 1580 33033
rect 130 32988 138 33022
rect 1572 32988 1580 33022
rect 130 32977 1580 32988
rect 130 32936 1580 32947
rect 130 32902 138 32936
rect 1572 32902 1580 32936
rect 130 32891 1580 32902
rect 130 32850 1580 32861
rect 130 32816 138 32850
rect 1572 32816 1580 32850
rect 130 32805 1580 32816
rect 130 32764 1580 32775
rect 130 32730 138 32764
rect 1572 32730 1580 32764
rect 130 32719 1580 32730
rect 130 32678 1580 32689
rect 130 32644 138 32678
rect 1572 32644 1580 32678
rect 130 32633 1580 32644
rect 130 32592 1580 32603
rect 130 32558 138 32592
rect 1572 32558 1580 32592
rect 130 32547 1580 32558
rect 130 32506 1580 32517
rect 130 32472 138 32506
rect 1572 32472 1580 32506
rect 130 32461 1580 32472
rect 130 32420 1580 32431
rect 130 32386 138 32420
rect 1572 32386 1580 32420
rect 130 32375 1580 32386
rect 130 32334 1580 32345
rect 130 32300 138 32334
rect 1572 32300 1580 32334
rect 130 32289 1580 32300
rect 130 32248 1580 32259
rect 130 32214 138 32248
rect 1572 32214 1580 32248
rect 130 32203 1580 32214
rect 130 32162 1580 32173
rect 130 32128 138 32162
rect 1572 32128 1580 32162
rect 130 32117 1580 32128
rect 130 32076 1580 32087
rect 130 32042 138 32076
rect 1572 32042 1580 32076
rect 130 32031 1580 32042
rect 130 31990 1580 32001
rect 130 31956 138 31990
rect 1572 31956 1580 31990
rect 130 31945 1580 31956
rect 130 31904 1580 31915
rect 130 31870 138 31904
rect 1572 31870 1580 31904
rect 130 31859 1580 31870
rect 130 31818 1580 31829
rect 130 31784 138 31818
rect 1572 31784 1580 31818
rect 130 31773 1580 31784
rect 130 31732 1580 31743
rect 130 31698 138 31732
rect 1572 31698 1580 31732
rect 130 31687 1580 31698
rect 130 31646 1580 31657
rect 130 31612 138 31646
rect 1572 31612 1580 31646
rect 130 31601 1580 31612
rect 130 31560 1580 31571
rect 130 31526 138 31560
rect 1572 31526 1580 31560
rect 130 31515 1580 31526
rect 130 31474 1580 31485
rect 130 31440 138 31474
rect 1572 31440 1580 31474
rect 130 31429 1580 31440
rect 130 31388 1580 31399
rect 130 31354 138 31388
rect 1572 31354 1580 31388
rect 130 31343 1580 31354
rect 130 31302 1580 31313
rect 130 31268 138 31302
rect 1572 31268 1580 31302
rect 130 31257 1580 31268
rect 130 31216 1580 31227
rect 130 31182 138 31216
rect 1572 31182 1580 31216
rect 130 31171 1580 31182
rect 130 31130 1580 31141
rect 130 31096 138 31130
rect 1572 31096 1580 31130
rect 130 31085 1580 31096
rect 130 31044 1580 31055
rect 130 31010 138 31044
rect 1572 31010 1580 31044
rect 130 30999 1580 31010
rect 130 30958 1580 30969
rect 130 30924 138 30958
rect 1572 30924 1580 30958
rect 130 30913 1580 30924
rect 130 30872 1580 30883
rect 130 30838 138 30872
rect 1572 30838 1580 30872
rect 130 30827 1580 30838
rect 130 30786 1580 30797
rect 130 30752 138 30786
rect 1572 30752 1580 30786
rect 130 30741 1580 30752
rect 130 30700 1580 30711
rect 130 30666 138 30700
rect 1572 30666 1580 30700
rect 130 30655 1580 30666
rect 130 30614 1580 30625
rect 130 30580 138 30614
rect 1572 30580 1580 30614
rect 130 30569 1580 30580
rect 130 30528 1580 30539
rect 130 30494 138 30528
rect 1572 30494 1580 30528
rect 130 30483 1580 30494
rect 130 30442 1580 30453
rect 130 30408 138 30442
rect 1572 30408 1580 30442
rect 130 30397 1580 30408
rect 130 30356 1580 30367
rect 130 30322 138 30356
rect 1572 30322 1580 30356
rect 130 30311 1580 30322
rect 130 30270 1580 30281
rect 130 30236 138 30270
rect 1572 30236 1580 30270
rect 130 30225 1580 30236
rect 130 30184 1580 30195
rect 130 30150 138 30184
rect 1572 30150 1580 30184
rect 130 30139 1580 30150
rect 130 30098 1580 30109
rect 130 30064 138 30098
rect 1572 30064 1580 30098
rect 130 30053 1580 30064
rect 130 30012 1580 30023
rect 130 29978 138 30012
rect 1572 29978 1580 30012
rect 130 29967 1580 29978
rect 130 29926 1580 29937
rect 130 29892 138 29926
rect 1572 29892 1580 29926
rect 130 29881 1580 29892
rect 130 29840 1580 29851
rect 130 29806 138 29840
rect 1572 29806 1580 29840
rect 130 29795 1580 29806
rect 130 29754 1580 29765
rect 130 29720 138 29754
rect 1572 29720 1580 29754
rect 130 29709 1580 29720
rect 130 29668 1580 29679
rect 130 29634 138 29668
rect 1572 29634 1580 29668
rect 130 29623 1580 29634
rect 130 29582 1580 29593
rect 130 29548 138 29582
rect 1572 29548 1580 29582
rect 130 29537 1580 29548
rect 130 29496 1580 29507
rect 130 29462 138 29496
rect 1572 29462 1580 29496
rect 130 29451 1580 29462
rect 130 29410 1580 29421
rect 130 29376 138 29410
rect 1572 29376 1580 29410
rect 130 29365 1580 29376
rect 130 29324 1580 29335
rect 130 29290 138 29324
rect 1572 29290 1580 29324
rect 130 29279 1580 29290
rect 130 29238 1580 29249
rect 130 29204 138 29238
rect 1572 29204 1580 29238
rect 130 29193 1580 29204
rect 130 29152 1580 29163
rect 130 29118 138 29152
rect 1572 29118 1580 29152
rect 130 29107 1580 29118
rect 130 29066 1580 29077
rect 130 29032 138 29066
rect 1572 29032 1580 29066
rect 130 29021 1580 29032
rect 130 28980 1580 28991
rect 130 28946 138 28980
rect 1572 28946 1580 28980
rect 130 28935 1580 28946
rect 130 28894 1580 28905
rect 130 28860 138 28894
rect 1572 28860 1580 28894
rect 130 28849 1580 28860
rect 130 28808 1580 28819
rect 130 28774 138 28808
rect 1572 28774 1580 28808
rect 130 28763 1580 28774
rect 130 28722 1580 28733
rect 130 28688 138 28722
rect 1572 28688 1580 28722
rect 130 28677 1580 28688
rect 130 28636 1580 28647
rect 130 28602 138 28636
rect 1572 28602 1580 28636
rect 130 28591 1580 28602
rect 130 28550 1580 28561
rect 130 28516 138 28550
rect 1572 28516 1580 28550
rect 130 28505 1580 28516
rect 130 28464 1580 28475
rect 130 28430 138 28464
rect 1572 28430 1580 28464
rect 130 28419 1580 28430
rect 130 28378 1580 28389
rect 130 28344 138 28378
rect 1572 28344 1580 28378
rect 130 28333 1580 28344
rect 130 28292 1580 28303
rect 130 28258 138 28292
rect 1572 28258 1580 28292
rect 130 28247 1580 28258
rect 130 28206 1580 28217
rect 130 28172 138 28206
rect 1572 28172 1580 28206
rect 130 28161 1580 28172
rect 130 28120 1580 28131
rect 130 28086 138 28120
rect 1572 28086 1580 28120
rect 130 28075 1580 28086
rect 130 28034 1580 28045
rect 130 28000 138 28034
rect 1572 28000 1580 28034
rect 130 27989 1580 28000
rect 130 27948 1580 27959
rect 130 27914 138 27948
rect 1572 27914 1580 27948
rect 130 27903 1580 27914
rect 130 27862 1580 27873
rect 130 27828 138 27862
rect 1572 27828 1580 27862
rect 130 27817 1580 27828
rect 130 27776 1580 27787
rect 130 27742 138 27776
rect 1572 27742 1580 27776
rect 130 27731 1580 27742
rect 130 27690 1580 27701
rect 130 27656 138 27690
rect 1572 27656 1580 27690
rect 130 27645 1580 27656
rect 130 27604 1580 27615
rect 130 27570 138 27604
rect 1572 27570 1580 27604
rect 130 27559 1580 27570
rect 130 27518 1580 27529
rect 130 27484 138 27518
rect 1572 27484 1580 27518
rect 130 27473 1580 27484
rect 130 27432 1580 27443
rect 130 27398 138 27432
rect 1572 27398 1580 27432
rect 130 27387 1580 27398
rect 130 27346 1580 27357
rect 130 27312 138 27346
rect 1572 27312 1580 27346
rect 130 27301 1580 27312
rect 130 27260 1580 27271
rect 130 27226 138 27260
rect 1572 27226 1580 27260
rect 130 27215 1580 27226
rect 130 27174 1580 27185
rect 130 27140 138 27174
rect 1572 27140 1580 27174
rect 130 27129 1580 27140
rect 130 27088 1580 27099
rect 130 27054 138 27088
rect 1572 27054 1580 27088
rect 130 27043 1580 27054
rect 130 27002 1580 27013
rect 130 26968 138 27002
rect 1572 26968 1580 27002
rect 130 26957 1580 26968
rect 130 26916 1580 26927
rect 130 26882 138 26916
rect 1572 26882 1580 26916
rect 130 26871 1580 26882
rect 130 26830 1580 26841
rect 130 26796 138 26830
rect 1572 26796 1580 26830
rect 130 26785 1580 26796
rect 130 26744 1580 26755
rect 130 26710 138 26744
rect 1572 26710 1580 26744
rect 130 26699 1580 26710
rect 130 26658 1580 26669
rect 130 26624 138 26658
rect 1572 26624 1580 26658
rect 130 26613 1580 26624
rect 130 26572 1580 26583
rect 130 26538 138 26572
rect 1572 26538 1580 26572
rect 130 26527 1580 26538
rect 130 26486 1580 26497
rect 130 26452 138 26486
rect 1572 26452 1580 26486
rect 130 26441 1580 26452
rect 130 26400 1580 26411
rect 130 26366 138 26400
rect 1572 26366 1580 26400
rect 130 26355 1580 26366
rect 130 26314 1580 26325
rect 130 26280 138 26314
rect 1572 26280 1580 26314
rect 130 26269 1580 26280
rect 130 26228 1580 26239
rect 130 26194 138 26228
rect 1572 26194 1580 26228
rect 130 26183 1580 26194
rect 130 26142 1580 26153
rect 130 26108 138 26142
rect 1572 26108 1580 26142
rect 130 26097 1580 26108
rect 130 26056 1580 26067
rect 130 26022 138 26056
rect 1572 26022 1580 26056
rect 130 26011 1580 26022
rect 130 25970 1580 25981
rect 130 25936 138 25970
rect 1572 25936 1580 25970
rect 130 25925 1580 25936
rect 130 25884 1580 25895
rect 130 25850 138 25884
rect 1572 25850 1580 25884
rect 130 25839 1580 25850
rect 130 25798 1580 25809
rect 130 25764 138 25798
rect 1572 25764 1580 25798
rect 130 25753 1580 25764
rect 130 25712 1580 25723
rect 130 25678 138 25712
rect 1572 25678 1580 25712
rect 130 25667 1580 25678
rect 130 25626 1580 25637
rect 130 25592 138 25626
rect 1572 25592 1580 25626
rect 130 25581 1580 25592
rect 130 25540 1580 25551
rect 130 25506 138 25540
rect 1572 25506 1580 25540
rect 130 25495 1580 25506
rect 130 25454 1580 25465
rect 130 25420 138 25454
rect 1572 25420 1580 25454
rect 130 25409 1580 25420
rect 130 25368 1580 25379
rect 130 25334 138 25368
rect 1572 25334 1580 25368
rect 130 25323 1580 25334
rect 130 25282 1580 25293
rect 130 25248 138 25282
rect 1572 25248 1580 25282
rect 130 25237 1580 25248
rect 130 25196 1580 25207
rect 130 25162 138 25196
rect 1572 25162 1580 25196
rect 130 25151 1580 25162
rect 130 25110 1580 25121
rect 130 25076 138 25110
rect 1572 25076 1580 25110
rect 130 25065 1580 25076
rect 130 25024 1580 25035
rect 130 24990 138 25024
rect 1572 24990 1580 25024
rect 130 24979 1580 24990
rect 130 24938 1580 24949
rect 130 24904 138 24938
rect 1572 24904 1580 24938
rect 130 24893 1580 24904
rect 130 24852 1580 24863
rect 130 24818 138 24852
rect 1572 24818 1580 24852
rect 130 24807 1580 24818
rect 130 24766 1580 24777
rect 130 24732 138 24766
rect 1572 24732 1580 24766
rect 130 24721 1580 24732
rect 130 24680 1580 24691
rect 130 24646 138 24680
rect 1572 24646 1580 24680
rect 130 24635 1580 24646
rect 130 24594 1580 24605
rect 130 24560 138 24594
rect 1572 24560 1580 24594
rect 130 24549 1580 24560
rect 130 24508 1580 24519
rect 130 24474 138 24508
rect 1572 24474 1580 24508
rect 130 24463 1580 24474
rect 130 24422 1580 24433
rect 130 24388 138 24422
rect 1572 24388 1580 24422
rect 130 24377 1580 24388
rect 130 24336 1580 24347
rect 130 24302 138 24336
rect 1572 24302 1580 24336
rect 130 24291 1580 24302
rect 130 24250 1580 24261
rect 130 24216 138 24250
rect 1572 24216 1580 24250
rect 130 24205 1580 24216
rect 130 24164 1580 24175
rect 130 24130 138 24164
rect 1572 24130 1580 24164
rect 130 24119 1580 24130
rect 130 24078 1580 24089
rect 130 24044 138 24078
rect 1572 24044 1580 24078
rect 130 24033 1580 24044
rect 130 23992 1580 24003
rect 130 23958 138 23992
rect 1572 23958 1580 23992
rect 130 23947 1580 23958
rect 130 23906 1580 23917
rect 130 23872 138 23906
rect 1572 23872 1580 23906
rect 130 23861 1580 23872
rect 130 23820 1580 23831
rect 130 23786 138 23820
rect 1572 23786 1580 23820
rect 130 23775 1580 23786
rect 130 23734 1580 23745
rect 130 23700 138 23734
rect 1572 23700 1580 23734
rect 130 23689 1580 23700
rect 130 23648 1580 23659
rect 130 23614 138 23648
rect 1572 23614 1580 23648
rect 130 23603 1580 23614
rect 130 23562 1580 23573
rect 130 23528 138 23562
rect 1572 23528 1580 23562
rect 130 23517 1580 23528
rect 130 23476 1580 23487
rect 130 23442 138 23476
rect 1572 23442 1580 23476
rect 130 23431 1580 23442
rect 130 23390 1580 23401
rect 130 23356 138 23390
rect 1572 23356 1580 23390
rect 130 23345 1580 23356
rect 130 23304 1580 23315
rect 130 23270 138 23304
rect 1572 23270 1580 23304
rect 130 23259 1580 23270
rect 130 23218 1580 23229
rect 130 23184 138 23218
rect 1572 23184 1580 23218
rect 130 23173 1580 23184
rect 130 23132 1580 23143
rect 130 23098 138 23132
rect 1572 23098 1580 23132
rect 130 23087 1580 23098
rect 130 23046 1580 23057
rect 130 23012 138 23046
rect 1572 23012 1580 23046
rect 130 23001 1580 23012
rect 130 22960 1580 22971
rect 130 22926 138 22960
rect 1572 22926 1580 22960
rect 130 22915 1580 22926
rect 130 22874 1580 22885
rect 130 22840 138 22874
rect 1572 22840 1580 22874
rect 130 22829 1580 22840
rect 130 22788 1580 22799
rect 130 22754 138 22788
rect 1572 22754 1580 22788
rect 130 22743 1580 22754
rect 130 22702 1580 22713
rect 130 22668 138 22702
rect 1572 22668 1580 22702
rect 130 22657 1580 22668
rect 130 22616 1580 22627
rect 130 22582 138 22616
rect 1572 22582 1580 22616
rect 130 22571 1580 22582
rect 130 22530 1580 22541
rect 130 22496 138 22530
rect 1572 22496 1580 22530
rect 130 22485 1580 22496
rect 130 22444 1580 22455
rect 130 22410 138 22444
rect 1572 22410 1580 22444
rect 130 22399 1580 22410
rect 130 22358 1580 22369
rect 130 22324 138 22358
rect 1572 22324 1580 22358
rect 130 22313 1580 22324
rect 130 22272 1580 22283
rect 130 22238 138 22272
rect 1572 22238 1580 22272
rect 130 22227 1580 22238
rect 130 22186 1580 22197
rect 130 22152 138 22186
rect 1572 22152 1580 22186
rect 130 22141 1580 22152
rect 130 22100 1580 22111
rect 130 22066 138 22100
rect 1572 22066 1580 22100
rect 130 22055 1580 22066
rect 130 22014 1580 22025
rect 130 21980 138 22014
rect 1572 21980 1580 22014
rect 130 21969 1580 21980
rect 130 21928 1580 21939
rect 130 21894 138 21928
rect 1572 21894 1580 21928
rect 130 21883 1580 21894
rect 130 21842 1580 21853
rect 130 21808 138 21842
rect 1572 21808 1580 21842
rect 130 21797 1580 21808
rect 130 21756 1580 21767
rect 130 21722 138 21756
rect 1572 21722 1580 21756
rect 130 21711 1580 21722
rect 130 21670 1580 21681
rect 130 21636 138 21670
rect 1572 21636 1580 21670
rect 130 21625 1580 21636
rect 130 21584 1580 21595
rect 130 21550 138 21584
rect 1572 21550 1580 21584
rect 130 21539 1580 21550
rect 130 21498 1580 21509
rect 130 21464 138 21498
rect 1572 21464 1580 21498
rect 130 21453 1580 21464
rect 130 21412 1580 21423
rect 130 21378 138 21412
rect 1572 21378 1580 21412
rect 130 21367 1580 21378
rect 130 21326 1580 21337
rect 130 21292 138 21326
rect 1572 21292 1580 21326
rect 130 21281 1580 21292
rect 130 21240 1580 21251
rect 130 21206 138 21240
rect 1572 21206 1580 21240
rect 130 21195 1580 21206
rect 130 21154 1580 21165
rect 130 21120 138 21154
rect 1572 21120 1580 21154
rect 130 21109 1580 21120
rect 130 21068 1580 21079
rect 130 21034 138 21068
rect 1572 21034 1580 21068
rect 130 21023 1580 21034
rect 130 20982 1580 20993
rect 130 20948 138 20982
rect 1572 20948 1580 20982
rect 130 20937 1580 20948
rect 130 20896 1580 20907
rect 130 20862 138 20896
rect 1572 20862 1580 20896
rect 130 20851 1580 20862
rect 130 20810 1580 20821
rect 130 20776 138 20810
rect 1572 20776 1580 20810
rect 130 20765 1580 20776
rect 130 20724 1580 20735
rect 130 20690 138 20724
rect 1572 20690 1580 20724
rect 130 20679 1580 20690
rect 130 20638 1580 20649
rect 130 20604 138 20638
rect 1572 20604 1580 20638
rect 130 20593 1580 20604
rect 130 20552 1580 20563
rect 130 20518 138 20552
rect 1572 20518 1580 20552
rect 130 20507 1580 20518
rect 130 20466 1580 20477
rect 130 20432 138 20466
rect 1572 20432 1580 20466
rect 130 20421 1580 20432
rect 130 20380 1580 20391
rect 130 20346 138 20380
rect 1572 20346 1580 20380
rect 130 20335 1580 20346
rect 130 20294 1580 20305
rect 130 20260 138 20294
rect 1572 20260 1580 20294
rect 130 20249 1580 20260
rect 130 20208 1580 20219
rect 130 20174 138 20208
rect 1572 20174 1580 20208
rect 130 20163 1580 20174
rect 130 20122 1580 20133
rect 130 20088 138 20122
rect 1572 20088 1580 20122
rect 130 20077 1580 20088
rect 130 20036 1580 20047
rect 130 20002 138 20036
rect 1572 20002 1580 20036
rect 130 19991 1580 20002
rect 130 19950 1580 19961
rect 130 19916 138 19950
rect 1572 19916 1580 19950
rect 130 19905 1580 19916
rect 130 19864 1580 19875
rect 130 19830 138 19864
rect 1572 19830 1580 19864
rect 130 19819 1580 19830
rect 130 19778 1580 19789
rect 130 19744 138 19778
rect 1572 19744 1580 19778
rect 130 19733 1580 19744
rect 130 19692 1580 19703
rect 130 19658 138 19692
rect 1572 19658 1580 19692
rect 130 19647 1580 19658
rect 130 19606 1580 19617
rect 130 19572 138 19606
rect 1572 19572 1580 19606
rect 130 19561 1580 19572
rect 130 19520 1580 19531
rect 130 19486 138 19520
rect 1572 19486 1580 19520
rect 130 19475 1580 19486
rect 130 19434 1580 19445
rect 130 19400 138 19434
rect 1572 19400 1580 19434
rect 130 19389 1580 19400
rect 130 19348 1580 19359
rect 130 19314 138 19348
rect 1572 19314 1580 19348
rect 130 19303 1580 19314
rect 130 19262 1580 19273
rect 130 19228 138 19262
rect 1572 19228 1580 19262
rect 130 19217 1580 19228
rect 130 19176 1580 19187
rect 130 19142 138 19176
rect 1572 19142 1580 19176
rect 130 19131 1580 19142
rect 130 19090 1580 19101
rect 130 19056 138 19090
rect 1572 19056 1580 19090
rect 130 19045 1580 19056
rect 130 19004 1580 19015
rect 130 18970 138 19004
rect 1572 18970 1580 19004
rect 130 18959 1580 18970
rect 130 18918 1580 18929
rect 130 18884 138 18918
rect 1572 18884 1580 18918
rect 130 18873 1580 18884
rect 130 18832 1580 18843
rect 130 18798 138 18832
rect 1572 18798 1580 18832
rect 130 18787 1580 18798
rect 130 18746 1580 18757
rect 130 18712 138 18746
rect 1572 18712 1580 18746
rect 130 18701 1580 18712
rect 130 18660 1580 18671
rect 130 18626 138 18660
rect 1572 18626 1580 18660
rect 130 18615 1580 18626
rect 130 18574 1580 18585
rect 130 18540 138 18574
rect 1572 18540 1580 18574
rect 130 18529 1580 18540
rect 130 18488 1580 18499
rect 130 18454 138 18488
rect 1572 18454 1580 18488
rect 130 18443 1580 18454
rect 130 18402 1580 18413
rect 130 18368 138 18402
rect 1572 18368 1580 18402
rect 130 18357 1580 18368
rect 130 18316 1580 18327
rect 130 18282 138 18316
rect 1572 18282 1580 18316
rect 130 18271 1580 18282
rect 130 18230 1580 18241
rect 130 18196 138 18230
rect 1572 18196 1580 18230
rect 130 18185 1580 18196
rect 130 18144 1580 18155
rect 130 18110 138 18144
rect 1572 18110 1580 18144
rect 130 18099 1580 18110
rect 130 18058 1580 18069
rect 130 18024 138 18058
rect 1572 18024 1580 18058
rect 130 18013 1580 18024
rect 130 17972 1580 17983
rect 130 17938 138 17972
rect 1572 17938 1580 17972
rect 130 17927 1580 17938
rect 130 17886 1580 17897
rect 130 17852 138 17886
rect 1572 17852 1580 17886
rect 130 17841 1580 17852
rect 130 17800 1580 17811
rect 130 17766 138 17800
rect 1572 17766 1580 17800
rect 130 17755 1580 17766
rect 130 17714 1580 17725
rect 130 17680 138 17714
rect 1572 17680 1580 17714
rect 130 17669 1580 17680
rect 130 17628 1580 17639
rect 130 17594 138 17628
rect 1572 17594 1580 17628
rect 130 17583 1580 17594
rect 130 17542 1580 17553
rect 130 17508 138 17542
rect 1572 17508 1580 17542
rect 130 17497 1580 17508
rect 130 17456 1580 17467
rect 130 17422 138 17456
rect 1572 17422 1580 17456
rect 130 17411 1580 17422
rect 130 17370 1580 17381
rect 130 17336 138 17370
rect 1572 17336 1580 17370
rect 130 17325 1580 17336
rect 130 17284 1580 17295
rect 130 17250 138 17284
rect 1572 17250 1580 17284
rect 130 17239 1580 17250
rect 130 17198 1580 17209
rect 130 17164 138 17198
rect 1572 17164 1580 17198
rect 130 17153 1580 17164
rect 130 17112 1580 17123
rect 130 17078 138 17112
rect 1572 17078 1580 17112
rect 130 17067 1580 17078
rect 130 17026 1580 17037
rect 130 16992 138 17026
rect 1572 16992 1580 17026
rect 130 16981 1580 16992
rect 130 16940 1580 16951
rect 130 16906 138 16940
rect 1572 16906 1580 16940
rect 130 16895 1580 16906
rect 130 16854 1580 16865
rect 130 16820 138 16854
rect 1572 16820 1580 16854
rect 130 16809 1580 16820
rect 130 16768 1580 16779
rect 130 16734 138 16768
rect 1572 16734 1580 16768
rect 130 16723 1580 16734
rect 130 16682 1580 16693
rect 130 16648 138 16682
rect 1572 16648 1580 16682
rect 130 16637 1580 16648
rect 130 16596 1580 16607
rect 130 16562 138 16596
rect 1572 16562 1580 16596
rect 130 16551 1580 16562
rect 130 16510 1580 16521
rect 130 16476 138 16510
rect 1572 16476 1580 16510
rect 130 16465 1580 16476
rect 130 16424 1580 16435
rect 130 16390 138 16424
rect 1572 16390 1580 16424
rect 130 16379 1580 16390
rect 130 16338 1580 16349
rect 130 16304 138 16338
rect 1572 16304 1580 16338
rect 130 16293 1580 16304
rect 130 16252 1580 16263
rect 130 16218 138 16252
rect 1572 16218 1580 16252
rect 130 16207 1580 16218
rect 130 16166 1580 16177
rect 130 16132 138 16166
rect 1572 16132 1580 16166
rect 130 16121 1580 16132
rect 130 16080 1580 16091
rect 130 16046 138 16080
rect 1572 16046 1580 16080
rect 130 16035 1580 16046
rect 130 15994 1580 16005
rect 130 15960 138 15994
rect 1572 15960 1580 15994
rect 130 15949 1580 15960
rect 130 15908 1580 15919
rect 130 15874 138 15908
rect 1572 15874 1580 15908
rect 130 15863 1580 15874
rect 130 15822 1580 15833
rect 130 15788 138 15822
rect 1572 15788 1580 15822
rect 130 15777 1580 15788
rect 130 15736 1580 15747
rect 130 15702 138 15736
rect 1572 15702 1580 15736
rect 130 15691 1580 15702
rect 130 15650 1580 15661
rect 130 15616 138 15650
rect 1572 15616 1580 15650
rect 130 15605 1580 15616
rect 130 15564 1580 15575
rect 130 15530 138 15564
rect 1572 15530 1580 15564
rect 130 15519 1580 15530
rect 130 15478 1580 15489
rect 130 15444 138 15478
rect 1572 15444 1580 15478
rect 130 15433 1580 15444
rect 130 15392 1580 15403
rect 130 15358 138 15392
rect 1572 15358 1580 15392
rect 130 15347 1580 15358
rect 130 15306 1580 15317
rect 130 15272 138 15306
rect 1572 15272 1580 15306
rect 130 15261 1580 15272
rect 130 15220 1580 15231
rect 130 15186 138 15220
rect 1572 15186 1580 15220
rect 130 15175 1580 15186
rect 130 15134 1580 15145
rect 130 15100 138 15134
rect 1572 15100 1580 15134
rect 130 15089 1580 15100
rect 130 15048 1580 15059
rect 130 15014 138 15048
rect 1572 15014 1580 15048
rect 130 15003 1580 15014
rect 130 14962 1580 14973
rect 130 14928 138 14962
rect 1572 14928 1580 14962
rect 130 14917 1580 14928
rect 130 14876 1580 14887
rect 130 14842 138 14876
rect 1572 14842 1580 14876
rect 130 14831 1580 14842
rect 130 14790 1580 14801
rect 130 14756 138 14790
rect 1572 14756 1580 14790
rect 130 14745 1580 14756
rect 130 14704 1580 14715
rect 130 14670 138 14704
rect 1572 14670 1580 14704
rect 130 14659 1580 14670
rect 130 14618 1580 14629
rect 130 14584 138 14618
rect 1572 14584 1580 14618
rect 130 14573 1580 14584
rect 130 14532 1580 14543
rect 130 14498 138 14532
rect 1572 14498 1580 14532
rect 130 14487 1580 14498
rect 130 14446 1580 14457
rect 130 14412 138 14446
rect 1572 14412 1580 14446
rect 130 14401 1580 14412
rect 130 14360 1580 14371
rect 130 14326 138 14360
rect 1572 14326 1580 14360
rect 130 14315 1580 14326
rect 130 14274 1580 14285
rect 130 14240 138 14274
rect 1572 14240 1580 14274
rect 130 14229 1580 14240
rect 130 14188 1580 14199
rect 130 14154 138 14188
rect 1572 14154 1580 14188
rect 130 14143 1580 14154
rect 130 14102 1580 14113
rect 130 14068 138 14102
rect 1572 14068 1580 14102
rect 130 14057 1580 14068
rect 130 14016 1580 14027
rect 130 13982 138 14016
rect 1572 13982 1580 14016
rect 130 13971 1580 13982
rect 130 13930 1580 13941
rect 130 13896 138 13930
rect 1572 13896 1580 13930
rect 130 13885 1580 13896
rect 130 13844 1580 13855
rect 130 13810 138 13844
rect 1572 13810 1580 13844
rect 130 13799 1580 13810
rect 130 13758 1580 13769
rect 130 13724 138 13758
rect 1572 13724 1580 13758
rect 130 13713 1580 13724
rect 130 13672 1580 13683
rect 130 13638 138 13672
rect 1572 13638 1580 13672
rect 130 13627 1580 13638
rect 130 13586 1580 13597
rect 130 13552 138 13586
rect 1572 13552 1580 13586
rect 130 13541 1580 13552
rect 130 13500 1580 13511
rect 130 13466 138 13500
rect 1572 13466 1580 13500
rect 130 13455 1580 13466
rect 130 13414 1580 13425
rect 130 13380 138 13414
rect 1572 13380 1580 13414
rect 130 13369 1580 13380
rect 130 13328 1580 13339
rect 130 13294 138 13328
rect 1572 13294 1580 13328
rect 130 13283 1580 13294
rect 130 13242 1580 13253
rect 130 13208 138 13242
rect 1572 13208 1580 13242
rect 130 13197 1580 13208
rect 130 13156 1580 13167
rect 130 13122 138 13156
rect 1572 13122 1580 13156
rect 130 13111 1580 13122
rect 130 13070 1580 13081
rect 130 13036 138 13070
rect 1572 13036 1580 13070
rect 130 13025 1580 13036
rect 130 12984 1580 12995
rect 130 12950 138 12984
rect 1572 12950 1580 12984
rect 130 12939 1580 12950
rect 130 12898 1580 12909
rect 130 12864 138 12898
rect 1572 12864 1580 12898
rect 130 12853 1580 12864
rect 130 12812 1580 12823
rect 130 12778 138 12812
rect 1572 12778 1580 12812
rect 130 12767 1580 12778
rect 130 12726 1580 12737
rect 130 12692 138 12726
rect 1572 12692 1580 12726
rect 130 12681 1580 12692
rect 130 12640 1580 12651
rect 130 12606 138 12640
rect 1572 12606 1580 12640
rect 130 12595 1580 12606
rect 130 12554 1580 12565
rect 130 12520 138 12554
rect 1572 12520 1580 12554
rect 130 12509 1580 12520
rect 130 12468 1580 12479
rect 130 12434 138 12468
rect 1572 12434 1580 12468
rect 130 12423 1580 12434
rect 130 12382 1580 12393
rect 130 12348 138 12382
rect 1572 12348 1580 12382
rect 130 12337 1580 12348
rect 130 12296 1580 12307
rect 130 12262 138 12296
rect 1572 12262 1580 12296
rect 130 12251 1580 12262
rect 130 12210 1580 12221
rect 130 12176 138 12210
rect 1572 12176 1580 12210
rect 130 12165 1580 12176
rect 130 12124 1580 12135
rect 130 12090 138 12124
rect 1572 12090 1580 12124
rect 130 12079 1580 12090
rect 130 12038 1580 12049
rect 130 12004 138 12038
rect 1572 12004 1580 12038
rect 130 11993 1580 12004
rect 130 11952 1580 11963
rect 130 11918 138 11952
rect 1572 11918 1580 11952
rect 130 11907 1580 11918
rect 130 11866 1580 11877
rect 130 11832 138 11866
rect 1572 11832 1580 11866
rect 130 11821 1580 11832
rect 130 11780 1580 11791
rect 130 11746 138 11780
rect 1572 11746 1580 11780
rect 130 11735 1580 11746
rect 130 11694 1580 11705
rect 130 11660 138 11694
rect 1572 11660 1580 11694
rect 130 11649 1580 11660
rect 130 11608 1580 11619
rect 130 11574 138 11608
rect 1572 11574 1580 11608
rect 130 11563 1580 11574
rect 130 11522 1580 11533
rect 130 11488 138 11522
rect 1572 11488 1580 11522
rect 130 11477 1580 11488
rect 130 11436 1580 11447
rect 130 11402 138 11436
rect 1572 11402 1580 11436
rect 130 11391 1580 11402
rect 130 11350 1580 11361
rect 130 11316 138 11350
rect 1572 11316 1580 11350
rect 130 11305 1580 11316
rect 130 11264 1580 11275
rect 130 11230 138 11264
rect 1572 11230 1580 11264
rect 130 11219 1580 11230
rect 130 11178 1580 11189
rect 130 11144 138 11178
rect 1572 11144 1580 11178
rect 130 11133 1580 11144
rect 130 11092 1580 11103
rect 130 11058 138 11092
rect 1572 11058 1580 11092
rect 130 11047 1580 11058
rect 130 11006 1580 11017
rect 130 10972 138 11006
rect 1572 10972 1580 11006
rect 130 10961 1580 10972
rect 130 10920 1580 10931
rect 130 10886 138 10920
rect 1572 10886 1580 10920
rect 130 10875 1580 10886
rect 130 10834 1580 10845
rect 130 10800 138 10834
rect 1572 10800 1580 10834
rect 130 10789 1580 10800
rect 130 10748 1580 10759
rect 130 10714 138 10748
rect 1572 10714 1580 10748
rect 130 10703 1580 10714
rect 130 10662 1580 10673
rect 130 10628 138 10662
rect 1572 10628 1580 10662
rect 130 10617 1580 10628
rect 130 10576 1580 10587
rect 130 10542 138 10576
rect 1572 10542 1580 10576
rect 130 10531 1580 10542
rect 130 10490 1580 10501
rect 130 10456 138 10490
rect 1572 10456 1580 10490
rect 130 10445 1580 10456
rect 130 10404 1580 10415
rect 130 10370 138 10404
rect 1572 10370 1580 10404
rect 130 10359 1580 10370
rect 130 10318 1580 10329
rect 130 10284 138 10318
rect 1572 10284 1580 10318
rect 130 10273 1580 10284
rect 130 10232 1580 10243
rect 130 10198 138 10232
rect 1572 10198 1580 10232
rect 130 10187 1580 10198
rect 130 10146 1580 10157
rect 130 10112 138 10146
rect 1572 10112 1580 10146
rect 130 10101 1580 10112
rect 130 10060 1580 10071
rect 130 10026 138 10060
rect 1572 10026 1580 10060
rect 130 10015 1580 10026
rect 130 9974 1580 9985
rect 130 9940 138 9974
rect 1572 9940 1580 9974
rect 130 9929 1580 9940
rect 130 9888 1580 9899
rect 130 9854 138 9888
rect 1572 9854 1580 9888
rect 130 9843 1580 9854
rect 130 9802 1580 9813
rect 130 9768 138 9802
rect 1572 9768 1580 9802
rect 130 9757 1580 9768
rect 130 9716 1580 9727
rect 130 9682 138 9716
rect 1572 9682 1580 9716
rect 130 9671 1580 9682
rect 130 9630 1580 9641
rect 130 9596 138 9630
rect 1572 9596 1580 9630
rect 130 9585 1580 9596
rect 130 9544 1580 9555
rect 130 9510 138 9544
rect 1572 9510 1580 9544
rect 130 9499 1580 9510
rect 130 9458 1580 9469
rect 130 9424 138 9458
rect 1572 9424 1580 9458
rect 130 9413 1580 9424
rect 130 9372 1580 9383
rect 130 9338 138 9372
rect 1572 9338 1580 9372
rect 130 9327 1580 9338
rect 130 9286 1580 9297
rect 130 9252 138 9286
rect 1572 9252 1580 9286
rect 130 9241 1580 9252
rect 130 9200 1580 9211
rect 130 9166 138 9200
rect 1572 9166 1580 9200
rect 130 9155 1580 9166
rect 130 9114 1580 9125
rect 130 9080 138 9114
rect 1572 9080 1580 9114
rect 130 9069 1580 9080
rect 130 9028 1580 9039
rect 130 8994 138 9028
rect 1572 8994 1580 9028
rect 130 8983 1580 8994
rect 130 8942 1580 8953
rect 130 8908 138 8942
rect 1572 8908 1580 8942
rect 130 8897 1580 8908
rect 130 8856 1580 8867
rect 130 8822 138 8856
rect 1572 8822 1580 8856
rect 130 8811 1580 8822
rect 130 8770 1580 8781
rect 130 8736 138 8770
rect 1572 8736 1580 8770
rect 130 8725 1580 8736
rect 130 8684 1580 8695
rect 130 8650 138 8684
rect 1572 8650 1580 8684
rect 130 8639 1580 8650
rect 130 8598 1580 8609
rect 130 8564 138 8598
rect 1572 8564 1580 8598
rect 130 8553 1580 8564
rect 130 8512 1580 8523
rect 130 8478 138 8512
rect 1572 8478 1580 8512
rect 130 8467 1580 8478
rect 130 8426 1580 8437
rect 130 8392 138 8426
rect 1572 8392 1580 8426
rect 130 8381 1580 8392
rect 130 8340 1580 8351
rect 130 8306 138 8340
rect 1572 8306 1580 8340
rect 130 8295 1580 8306
rect 130 8254 1580 8265
rect 130 8220 138 8254
rect 1572 8220 1580 8254
rect 130 8209 1580 8220
rect 130 8168 1580 8179
rect 130 8134 138 8168
rect 1572 8134 1580 8168
rect 130 8123 1580 8134
rect 130 8082 1580 8093
rect 130 8048 138 8082
rect 1572 8048 1580 8082
rect 130 8037 1580 8048
rect 130 7996 1580 8007
rect 130 7962 138 7996
rect 1572 7962 1580 7996
rect 130 7951 1580 7962
rect 130 7910 1580 7921
rect 130 7876 138 7910
rect 1572 7876 1580 7910
rect 130 7865 1580 7876
rect 130 7824 1580 7835
rect 130 7790 138 7824
rect 1572 7790 1580 7824
rect 130 7779 1580 7790
rect 130 7738 1580 7749
rect 130 7704 138 7738
rect 1572 7704 1580 7738
rect 130 7693 1580 7704
rect 130 7652 1580 7663
rect 130 7618 138 7652
rect 1572 7618 1580 7652
rect 130 7607 1580 7618
rect 130 7566 1580 7577
rect 130 7532 138 7566
rect 1572 7532 1580 7566
rect 130 7521 1580 7532
rect 130 7480 1580 7491
rect 130 7446 138 7480
rect 1572 7446 1580 7480
rect 130 7435 1580 7446
rect 130 7394 1580 7405
rect 130 7360 138 7394
rect 1572 7360 1580 7394
rect 130 7349 1580 7360
rect 130 7308 1580 7319
rect 130 7274 138 7308
rect 1572 7274 1580 7308
rect 130 7263 1580 7274
rect 130 7222 1580 7233
rect 130 7188 138 7222
rect 1572 7188 1580 7222
rect 130 7177 1580 7188
rect 130 7136 1580 7147
rect 130 7102 138 7136
rect 1572 7102 1580 7136
rect 130 7091 1580 7102
rect 130 7050 1580 7061
rect 130 7016 138 7050
rect 1572 7016 1580 7050
rect 130 7005 1580 7016
rect 130 6964 1580 6975
rect 130 6930 138 6964
rect 1572 6930 1580 6964
rect 130 6919 1580 6930
rect 130 6878 1580 6889
rect 130 6844 138 6878
rect 1572 6844 1580 6878
rect 130 6833 1580 6844
rect 130 6792 1580 6803
rect 130 6758 138 6792
rect 1572 6758 1580 6792
rect 130 6747 1580 6758
rect 130 6706 1580 6717
rect 130 6672 138 6706
rect 1572 6672 1580 6706
rect 130 6661 1580 6672
rect 130 6620 1580 6631
rect 130 6586 138 6620
rect 1572 6586 1580 6620
rect 130 6575 1580 6586
rect 130 6534 1580 6545
rect 130 6500 138 6534
rect 1572 6500 1580 6534
rect 130 6489 1580 6500
rect 130 6448 1580 6459
rect 130 6414 138 6448
rect 1572 6414 1580 6448
rect 130 6403 1580 6414
rect 130 6362 1580 6373
rect 130 6328 138 6362
rect 1572 6328 1580 6362
rect 130 6317 1580 6328
rect 130 6276 1580 6287
rect 130 6242 138 6276
rect 1572 6242 1580 6276
rect 130 6231 1580 6242
rect 130 6190 1580 6201
rect 130 6156 138 6190
rect 1572 6156 1580 6190
rect 130 6145 1580 6156
rect 130 6104 1580 6115
rect 130 6070 138 6104
rect 1572 6070 1580 6104
rect 130 6059 1580 6070
rect 130 6018 1580 6029
rect 130 5984 138 6018
rect 1572 5984 1580 6018
rect 130 5973 1580 5984
rect 130 5932 1580 5943
rect 130 5898 138 5932
rect 1572 5898 1580 5932
rect 130 5887 1580 5898
rect 130 5846 1580 5857
rect 130 5812 138 5846
rect 1572 5812 1580 5846
rect 130 5801 1580 5812
rect 130 5760 1580 5771
rect 130 5726 138 5760
rect 1572 5726 1580 5760
rect 130 5715 1580 5726
rect 130 5674 1580 5685
rect 130 5640 138 5674
rect 1572 5640 1580 5674
rect 130 5629 1580 5640
rect 130 5588 1580 5599
rect 130 5554 138 5588
rect 1572 5554 1580 5588
rect 130 5543 1580 5554
rect 130 5502 1580 5513
rect 130 5468 138 5502
rect 1572 5468 1580 5502
rect 130 5457 1580 5468
rect 130 5416 1580 5427
rect 130 5382 138 5416
rect 1572 5382 1580 5416
rect 130 5371 1580 5382
rect 130 5330 1580 5341
rect 130 5296 138 5330
rect 1572 5296 1580 5330
rect 130 5285 1580 5296
rect 130 5244 1580 5255
rect 130 5210 138 5244
rect 1572 5210 1580 5244
rect 130 5199 1580 5210
rect 130 5158 1580 5169
rect 130 5124 138 5158
rect 1572 5124 1580 5158
rect 130 5113 1580 5124
rect 130 5072 1580 5083
rect 130 5038 138 5072
rect 1572 5038 1580 5072
rect 130 5027 1580 5038
rect 130 4986 1580 4997
rect 130 4952 138 4986
rect 1572 4952 1580 4986
rect 130 4941 1580 4952
rect 130 4900 1580 4911
rect 130 4866 138 4900
rect 1572 4866 1580 4900
rect 130 4855 1580 4866
rect 130 4814 1580 4825
rect 130 4780 138 4814
rect 1572 4780 1580 4814
rect 130 4769 1580 4780
rect 130 4728 1580 4739
rect 130 4694 138 4728
rect 1572 4694 1580 4728
rect 130 4683 1580 4694
rect 130 4642 1580 4653
rect 130 4608 138 4642
rect 1572 4608 1580 4642
rect 130 4597 1580 4608
rect 130 4556 1580 4567
rect 130 4522 138 4556
rect 1572 4522 1580 4556
rect 130 4511 1580 4522
rect 130 4470 1580 4481
rect 130 4436 138 4470
rect 1572 4436 1580 4470
rect 130 4425 1580 4436
rect 130 4384 1580 4395
rect 130 4350 138 4384
rect 1572 4350 1580 4384
rect 130 4339 1580 4350
rect 130 4298 1580 4309
rect 130 4264 138 4298
rect 1572 4264 1580 4298
rect 130 4253 1580 4264
rect 130 4212 1580 4223
rect 130 4178 138 4212
rect 1572 4178 1580 4212
rect 130 4167 1580 4178
rect 130 4126 1580 4137
rect 130 4092 138 4126
rect 1572 4092 1580 4126
rect 130 4081 1580 4092
rect 130 4040 1580 4051
rect 130 4006 138 4040
rect 1572 4006 1580 4040
rect 130 3995 1580 4006
rect 130 3954 1580 3965
rect 130 3920 138 3954
rect 1572 3920 1580 3954
rect 130 3909 1580 3920
rect 130 3868 1580 3879
rect 130 3834 138 3868
rect 1572 3834 1580 3868
rect 130 3823 1580 3834
rect 130 3782 1580 3793
rect 130 3748 138 3782
rect 1572 3748 1580 3782
rect 130 3737 1580 3748
rect 130 3696 1580 3707
rect 130 3662 138 3696
rect 1572 3662 1580 3696
rect 130 3651 1580 3662
rect 130 3610 1580 3621
rect 130 3576 138 3610
rect 1572 3576 1580 3610
rect 130 3565 1580 3576
rect 130 3524 1580 3535
rect 130 3490 138 3524
rect 1572 3490 1580 3524
rect 130 3479 1580 3490
rect 130 3438 1580 3449
rect 130 3404 138 3438
rect 1572 3404 1580 3438
rect 130 3393 1580 3404
rect 130 3352 1580 3363
rect 130 3318 138 3352
rect 1572 3318 1580 3352
rect 130 3307 1580 3318
rect 130 3266 1580 3277
rect 130 3232 138 3266
rect 1572 3232 1580 3266
rect 130 3221 1580 3232
rect 130 3180 1580 3191
rect 130 3146 138 3180
rect 1572 3146 1580 3180
rect 130 3135 1580 3146
rect 130 3094 1580 3105
rect 130 3060 138 3094
rect 1572 3060 1580 3094
rect 130 3049 1580 3060
rect 130 3008 1580 3019
rect 130 2974 138 3008
rect 1572 2974 1580 3008
rect 130 2963 1580 2974
rect 130 2922 1580 2933
rect 130 2888 138 2922
rect 1572 2888 1580 2922
rect 130 2877 1580 2888
rect 130 2836 1580 2847
rect 130 2802 138 2836
rect 1572 2802 1580 2836
rect 130 2791 1580 2802
rect 130 2750 1580 2761
rect 130 2716 138 2750
rect 1572 2716 1580 2750
rect 130 2705 1580 2716
rect 130 2664 1580 2675
rect 130 2630 138 2664
rect 1572 2630 1580 2664
rect 130 2619 1580 2630
rect 130 2578 1580 2589
rect 130 2544 138 2578
rect 1572 2544 1580 2578
rect 130 2533 1580 2544
rect 130 2492 1580 2503
rect 130 2458 138 2492
rect 1572 2458 1580 2492
rect 130 2447 1580 2458
rect 130 2406 1580 2417
rect 130 2372 138 2406
rect 1572 2372 1580 2406
rect 130 2361 1580 2372
rect 130 2320 1580 2331
rect 130 2286 138 2320
rect 1572 2286 1580 2320
rect 130 2275 1580 2286
rect 130 2234 1580 2245
rect 130 2200 138 2234
rect 1572 2200 1580 2234
rect 130 2189 1580 2200
rect 130 2148 1580 2159
rect 130 2114 138 2148
rect 1572 2114 1580 2148
rect 130 2103 1580 2114
rect 130 2062 1580 2073
rect 130 2028 138 2062
rect 1572 2028 1580 2062
rect 130 2017 1580 2028
rect 130 1976 1580 1987
rect 130 1942 138 1976
rect 1572 1942 1580 1976
rect 130 1931 1580 1942
rect 130 1890 1580 1901
rect 130 1856 138 1890
rect 1572 1856 1580 1890
rect 130 1845 1580 1856
rect 130 1804 1580 1815
rect 130 1770 138 1804
rect 1572 1770 1580 1804
rect 130 1759 1580 1770
rect 130 1718 1580 1729
rect 130 1684 138 1718
rect 1572 1684 1580 1718
rect 130 1673 1580 1684
rect 130 1632 1580 1643
rect 130 1598 138 1632
rect 1572 1598 1580 1632
rect 130 1587 1580 1598
rect 130 1546 1580 1557
rect 130 1512 138 1546
rect 1572 1512 1580 1546
rect 130 1501 1580 1512
rect 130 1460 1580 1471
rect 130 1426 138 1460
rect 1572 1426 1580 1460
rect 130 1415 1580 1426
rect 130 1374 1580 1385
rect 130 1340 138 1374
rect 1572 1340 1580 1374
rect 130 1329 1580 1340
rect 130 1288 1580 1299
rect 130 1254 138 1288
rect 1572 1254 1580 1288
rect 130 1243 1580 1254
rect 130 1202 1580 1213
rect 130 1168 138 1202
rect 1572 1168 1580 1202
rect 130 1157 1580 1168
rect 130 1116 1580 1127
rect 130 1082 138 1116
rect 1572 1082 1580 1116
rect 130 1071 1580 1082
rect 130 1030 1580 1041
rect 130 996 138 1030
rect 1572 996 1580 1030
rect 130 985 1580 996
rect 130 944 1580 955
rect 130 910 138 944
rect 1572 910 1580 944
rect 130 899 1580 910
rect 130 858 1580 869
rect 130 824 138 858
rect 1572 824 1580 858
rect 130 813 1580 824
rect 130 772 1580 783
rect 130 738 138 772
rect 1572 738 1580 772
rect 130 727 1580 738
rect 130 686 1580 697
rect 130 652 138 686
rect 1572 652 1580 686
rect 130 641 1580 652
rect 130 600 1580 611
rect 130 566 138 600
rect 1572 566 1580 600
rect 130 555 1580 566
rect 130 514 1580 525
rect 130 480 138 514
rect 1572 480 1580 514
rect 130 469 1580 480
rect 130 428 1580 439
rect 130 394 138 428
rect 1572 394 1580 428
rect 130 383 1580 394
rect 130 342 1580 353
rect 130 308 138 342
rect 1572 308 1580 342
rect 130 297 1580 308
rect 130 256 1580 267
rect 130 222 138 256
rect 1572 222 1580 256
rect 130 211 1580 222
rect 130 170 1580 181
rect 130 136 138 170
rect 1572 136 1580 170
rect 130 124 1580 136
<< pdiffc >>
rect 138 100068 1572 100102
rect 138 99982 1572 100016
rect 138 99896 1572 99930
rect 138 99810 1572 99844
rect 138 99724 1572 99758
rect 138 99638 1572 99672
rect 138 99552 1572 99586
rect 138 99466 1572 99500
rect 138 99380 1572 99414
rect 138 99294 1572 99328
rect 138 99208 1572 99242
rect 138 99122 1572 99156
rect 138 99036 1572 99070
rect 138 98950 1572 98984
rect 138 98864 1572 98898
rect 138 98778 1572 98812
rect 138 98692 1572 98726
rect 138 98606 1572 98640
rect 138 98520 1572 98554
rect 138 98434 1572 98468
rect 138 98348 1572 98382
rect 138 98262 1572 98296
rect 138 98176 1572 98210
rect 138 98090 1572 98124
rect 138 98004 1572 98038
rect 138 97918 1572 97952
rect 138 97832 1572 97866
rect 138 97746 1572 97780
rect 138 97660 1572 97694
rect 138 97574 1572 97608
rect 138 97488 1572 97522
rect 138 97402 1572 97436
rect 138 97316 1572 97350
rect 138 97230 1572 97264
rect 138 97144 1572 97178
rect 138 97058 1572 97092
rect 138 96972 1572 97006
rect 138 96886 1572 96920
rect 138 96800 1572 96834
rect 138 96714 1572 96748
rect 138 96628 1572 96662
rect 138 96542 1572 96576
rect 138 96456 1572 96490
rect 138 96370 1572 96404
rect 138 96284 1572 96318
rect 138 96198 1572 96232
rect 138 96112 1572 96146
rect 138 96026 1572 96060
rect 138 95940 1572 95974
rect 138 95854 1572 95888
rect 138 95768 1572 95802
rect 138 95682 1572 95716
rect 138 95596 1572 95630
rect 138 95510 1572 95544
rect 138 95424 1572 95458
rect 138 95338 1572 95372
rect 138 95252 1572 95286
rect 138 95166 1572 95200
rect 138 95080 1572 95114
rect 138 94994 1572 95028
rect 138 94908 1572 94942
rect 138 94822 1572 94856
rect 138 94736 1572 94770
rect 138 94650 1572 94684
rect 138 94564 1572 94598
rect 138 94478 1572 94512
rect 138 94392 1572 94426
rect 138 94306 1572 94340
rect 138 94220 1572 94254
rect 138 94134 1572 94168
rect 138 94048 1572 94082
rect 138 93962 1572 93996
rect 138 93876 1572 93910
rect 138 93790 1572 93824
rect 138 93704 1572 93738
rect 138 93618 1572 93652
rect 138 93532 1572 93566
rect 138 93446 1572 93480
rect 138 93360 1572 93394
rect 138 93274 1572 93308
rect 138 93188 1572 93222
rect 138 93102 1572 93136
rect 138 93016 1572 93050
rect 138 92930 1572 92964
rect 138 92844 1572 92878
rect 138 92758 1572 92792
rect 138 92672 1572 92706
rect 138 92586 1572 92620
rect 138 92500 1572 92534
rect 138 92414 1572 92448
rect 138 92328 1572 92362
rect 138 92242 1572 92276
rect 138 92156 1572 92190
rect 138 92070 1572 92104
rect 138 91984 1572 92018
rect 138 91898 1572 91932
rect 138 91812 1572 91846
rect 138 91726 1572 91760
rect 138 91640 1572 91674
rect 138 91554 1572 91588
rect 138 91468 1572 91502
rect 138 91382 1572 91416
rect 138 91296 1572 91330
rect 138 91210 1572 91244
rect 138 91124 1572 91158
rect 138 91038 1572 91072
rect 138 90952 1572 90986
rect 138 90866 1572 90900
rect 138 90780 1572 90814
rect 138 90694 1572 90728
rect 138 90608 1572 90642
rect 138 90522 1572 90556
rect 138 90436 1572 90470
rect 138 90350 1572 90384
rect 138 90264 1572 90298
rect 138 90178 1572 90212
rect 138 90092 1572 90126
rect 138 90006 1572 90040
rect 138 89920 1572 89954
rect 138 89834 1572 89868
rect 138 89748 1572 89782
rect 138 89662 1572 89696
rect 138 89576 1572 89610
rect 138 89490 1572 89524
rect 138 89404 1572 89438
rect 138 89318 1572 89352
rect 138 89232 1572 89266
rect 138 89146 1572 89180
rect 138 89060 1572 89094
rect 138 88974 1572 89008
rect 138 88888 1572 88922
rect 138 88802 1572 88836
rect 138 88716 1572 88750
rect 138 88630 1572 88664
rect 138 88544 1572 88578
rect 138 88458 1572 88492
rect 138 88372 1572 88406
rect 138 88286 1572 88320
rect 138 88200 1572 88234
rect 138 88114 1572 88148
rect 138 88028 1572 88062
rect 138 87942 1572 87976
rect 138 87856 1572 87890
rect 138 87770 1572 87804
rect 138 87684 1572 87718
rect 138 87598 1572 87632
rect 138 87512 1572 87546
rect 138 87426 1572 87460
rect 138 87340 1572 87374
rect 138 87254 1572 87288
rect 138 87168 1572 87202
rect 138 87082 1572 87116
rect 138 86996 1572 87030
rect 138 86910 1572 86944
rect 138 86824 1572 86858
rect 138 86738 1572 86772
rect 138 86652 1572 86686
rect 138 86566 1572 86600
rect 138 86480 1572 86514
rect 138 86394 1572 86428
rect 138 86308 1572 86342
rect 138 86222 1572 86256
rect 138 86136 1572 86170
rect 138 86050 1572 86084
rect 138 85964 1572 85998
rect 138 85878 1572 85912
rect 138 85792 1572 85826
rect 138 85706 1572 85740
rect 138 85620 1572 85654
rect 138 85534 1572 85568
rect 138 85448 1572 85482
rect 138 85362 1572 85396
rect 138 85276 1572 85310
rect 138 85190 1572 85224
rect 138 85104 1572 85138
rect 138 85018 1572 85052
rect 138 84932 1572 84966
rect 138 84846 1572 84880
rect 138 84760 1572 84794
rect 138 84674 1572 84708
rect 138 84588 1572 84622
rect 138 84502 1572 84536
rect 138 84416 1572 84450
rect 138 84330 1572 84364
rect 138 84244 1572 84278
rect 138 84158 1572 84192
rect 138 84072 1572 84106
rect 138 83986 1572 84020
rect 138 83900 1572 83934
rect 138 83814 1572 83848
rect 138 83728 1572 83762
rect 138 83642 1572 83676
rect 138 83556 1572 83590
rect 138 83470 1572 83504
rect 138 83384 1572 83418
rect 138 83298 1572 83332
rect 138 83212 1572 83246
rect 138 83126 1572 83160
rect 138 83040 1572 83074
rect 138 82954 1572 82988
rect 138 82868 1572 82902
rect 138 82782 1572 82816
rect 138 82696 1572 82730
rect 138 82610 1572 82644
rect 138 82524 1572 82558
rect 138 82438 1572 82472
rect 138 82352 1572 82386
rect 138 82266 1572 82300
rect 138 82180 1572 82214
rect 138 82094 1572 82128
rect 138 82008 1572 82042
rect 138 81922 1572 81956
rect 138 81836 1572 81870
rect 138 81750 1572 81784
rect 138 81664 1572 81698
rect 138 81578 1572 81612
rect 138 81492 1572 81526
rect 138 81406 1572 81440
rect 138 81320 1572 81354
rect 138 81234 1572 81268
rect 138 81148 1572 81182
rect 138 81062 1572 81096
rect 138 80976 1572 81010
rect 138 80890 1572 80924
rect 138 80804 1572 80838
rect 138 80718 1572 80752
rect 138 80632 1572 80666
rect 138 80546 1572 80580
rect 138 80460 1572 80494
rect 138 80374 1572 80408
rect 138 80288 1572 80322
rect 138 80202 1572 80236
rect 138 80116 1572 80150
rect 138 80030 1572 80064
rect 138 79944 1572 79978
rect 138 79858 1572 79892
rect 138 79772 1572 79806
rect 138 79686 1572 79720
rect 138 79600 1572 79634
rect 138 79514 1572 79548
rect 138 79428 1572 79462
rect 138 79342 1572 79376
rect 138 79256 1572 79290
rect 138 79170 1572 79204
rect 138 79084 1572 79118
rect 138 78998 1572 79032
rect 138 78912 1572 78946
rect 138 78826 1572 78860
rect 138 78740 1572 78774
rect 138 78654 1572 78688
rect 138 78568 1572 78602
rect 138 78482 1572 78516
rect 138 78396 1572 78430
rect 138 78310 1572 78344
rect 138 78224 1572 78258
rect 138 78138 1572 78172
rect 138 78052 1572 78086
rect 138 77966 1572 78000
rect 138 77880 1572 77914
rect 138 77794 1572 77828
rect 138 77708 1572 77742
rect 138 77622 1572 77656
rect 138 77536 1572 77570
rect 138 77450 1572 77484
rect 138 77364 1572 77398
rect 138 77278 1572 77312
rect 138 77192 1572 77226
rect 138 77106 1572 77140
rect 138 77020 1572 77054
rect 138 76934 1572 76968
rect 138 76848 1572 76882
rect 138 76762 1572 76796
rect 138 76676 1572 76710
rect 138 76590 1572 76624
rect 138 76504 1572 76538
rect 138 76418 1572 76452
rect 138 76332 1572 76366
rect 138 76246 1572 76280
rect 138 76160 1572 76194
rect 138 76074 1572 76108
rect 138 75988 1572 76022
rect 138 75902 1572 75936
rect 138 75816 1572 75850
rect 138 75730 1572 75764
rect 138 75644 1572 75678
rect 138 75558 1572 75592
rect 138 75472 1572 75506
rect 138 75386 1572 75420
rect 138 75300 1572 75334
rect 138 75214 1572 75248
rect 138 75128 1572 75162
rect 138 75042 1572 75076
rect 138 74956 1572 74990
rect 138 74870 1572 74904
rect 138 74784 1572 74818
rect 138 74698 1572 74732
rect 138 74612 1572 74646
rect 138 74526 1572 74560
rect 138 74440 1572 74474
rect 138 74354 1572 74388
rect 138 74268 1572 74302
rect 138 74182 1572 74216
rect 138 74096 1572 74130
rect 138 74010 1572 74044
rect 138 73924 1572 73958
rect 138 73838 1572 73872
rect 138 73752 1572 73786
rect 138 73666 1572 73700
rect 138 73580 1572 73614
rect 138 73494 1572 73528
rect 138 73408 1572 73442
rect 138 73322 1572 73356
rect 138 73236 1572 73270
rect 138 73150 1572 73184
rect 138 73064 1572 73098
rect 138 72978 1572 73012
rect 138 72892 1572 72926
rect 138 72806 1572 72840
rect 138 72720 1572 72754
rect 138 72634 1572 72668
rect 138 72548 1572 72582
rect 138 72462 1572 72496
rect 138 72376 1572 72410
rect 138 72290 1572 72324
rect 138 72204 1572 72238
rect 138 72118 1572 72152
rect 138 72032 1572 72066
rect 138 71946 1572 71980
rect 138 71860 1572 71894
rect 138 71774 1572 71808
rect 138 71688 1572 71722
rect 138 71602 1572 71636
rect 138 71516 1572 71550
rect 138 71430 1572 71464
rect 138 71344 1572 71378
rect 138 71258 1572 71292
rect 138 71172 1572 71206
rect 138 71086 1572 71120
rect 138 71000 1572 71034
rect 138 70914 1572 70948
rect 138 70828 1572 70862
rect 138 70742 1572 70776
rect 138 70656 1572 70690
rect 138 70570 1572 70604
rect 138 70484 1572 70518
rect 138 70398 1572 70432
rect 138 70312 1572 70346
rect 138 70226 1572 70260
rect 138 70140 1572 70174
rect 138 70054 1572 70088
rect 138 69968 1572 70002
rect 138 69882 1572 69916
rect 138 69796 1572 69830
rect 138 69710 1572 69744
rect 138 69624 1572 69658
rect 138 69538 1572 69572
rect 138 69452 1572 69486
rect 138 69366 1572 69400
rect 138 69280 1572 69314
rect 138 69194 1572 69228
rect 138 69108 1572 69142
rect 138 69022 1572 69056
rect 138 68936 1572 68970
rect 138 68850 1572 68884
rect 138 68764 1572 68798
rect 138 68678 1572 68712
rect 138 68592 1572 68626
rect 138 68506 1572 68540
rect 138 68420 1572 68454
rect 138 68334 1572 68368
rect 138 68248 1572 68282
rect 138 68162 1572 68196
rect 138 68076 1572 68110
rect 138 67990 1572 68024
rect 138 67904 1572 67938
rect 138 67818 1572 67852
rect 138 67732 1572 67766
rect 138 67646 1572 67680
rect 138 67560 1572 67594
rect 138 67474 1572 67508
rect 138 67388 1572 67422
rect 138 67302 1572 67336
rect 138 67216 1572 67250
rect 138 67130 1572 67164
rect 138 67044 1572 67078
rect 138 66958 1572 66992
rect 138 66872 1572 66906
rect 138 66786 1572 66820
rect 138 66700 1572 66734
rect 138 66614 1572 66648
rect 138 66528 1572 66562
rect 138 66442 1572 66476
rect 138 66356 1572 66390
rect 138 66270 1572 66304
rect 138 66184 1572 66218
rect 138 66098 1572 66132
rect 138 66012 1572 66046
rect 138 65926 1572 65960
rect 138 65840 1572 65874
rect 138 65754 1572 65788
rect 138 65668 1572 65702
rect 138 65582 1572 65616
rect 138 65496 1572 65530
rect 138 65410 1572 65444
rect 138 65324 1572 65358
rect 138 65238 1572 65272
rect 138 65152 1572 65186
rect 138 65066 1572 65100
rect 138 64980 1572 65014
rect 138 64894 1572 64928
rect 138 64808 1572 64842
rect 138 64722 1572 64756
rect 138 64636 1572 64670
rect 138 64550 1572 64584
rect 138 64464 1572 64498
rect 138 64378 1572 64412
rect 138 64292 1572 64326
rect 138 64206 1572 64240
rect 138 64120 1572 64154
rect 138 64034 1572 64068
rect 138 63948 1572 63982
rect 138 63862 1572 63896
rect 138 63776 1572 63810
rect 138 63690 1572 63724
rect 138 63604 1572 63638
rect 138 63518 1572 63552
rect 138 63432 1572 63466
rect 138 63346 1572 63380
rect 138 63260 1572 63294
rect 138 63174 1572 63208
rect 138 63088 1572 63122
rect 138 63002 1572 63036
rect 138 62916 1572 62950
rect 138 62830 1572 62864
rect 138 62744 1572 62778
rect 138 62658 1572 62692
rect 138 62572 1572 62606
rect 138 62486 1572 62520
rect 138 62400 1572 62434
rect 138 62314 1572 62348
rect 138 62228 1572 62262
rect 138 62142 1572 62176
rect 138 62056 1572 62090
rect 138 61970 1572 62004
rect 138 61884 1572 61918
rect 138 61798 1572 61832
rect 138 61712 1572 61746
rect 138 61626 1572 61660
rect 138 61540 1572 61574
rect 138 61454 1572 61488
rect 138 61368 1572 61402
rect 138 61282 1572 61316
rect 138 61196 1572 61230
rect 138 61110 1572 61144
rect 138 61024 1572 61058
rect 138 60938 1572 60972
rect 138 60852 1572 60886
rect 138 60766 1572 60800
rect 138 60680 1572 60714
rect 138 60594 1572 60628
rect 138 60508 1572 60542
rect 138 60422 1572 60456
rect 138 60336 1572 60370
rect 138 60250 1572 60284
rect 138 60164 1572 60198
rect 138 60078 1572 60112
rect 138 59992 1572 60026
rect 138 59906 1572 59940
rect 138 59820 1572 59854
rect 138 59734 1572 59768
rect 138 59648 1572 59682
rect 138 59562 1572 59596
rect 138 59476 1572 59510
rect 138 59390 1572 59424
rect 138 59304 1572 59338
rect 138 59218 1572 59252
rect 138 59132 1572 59166
rect 138 59046 1572 59080
rect 138 58960 1572 58994
rect 138 58874 1572 58908
rect 138 58788 1572 58822
rect 138 58702 1572 58736
rect 138 58616 1572 58650
rect 138 58530 1572 58564
rect 138 58444 1572 58478
rect 138 58358 1572 58392
rect 138 58272 1572 58306
rect 138 58186 1572 58220
rect 138 58100 1572 58134
rect 138 58014 1572 58048
rect 138 57928 1572 57962
rect 138 57842 1572 57876
rect 138 57756 1572 57790
rect 138 57670 1572 57704
rect 138 57584 1572 57618
rect 138 57498 1572 57532
rect 138 57412 1572 57446
rect 138 57326 1572 57360
rect 138 57240 1572 57274
rect 138 57154 1572 57188
rect 138 57068 1572 57102
rect 138 56982 1572 57016
rect 138 56896 1572 56930
rect 138 56810 1572 56844
rect 138 56724 1572 56758
rect 138 56638 1572 56672
rect 138 56552 1572 56586
rect 138 56466 1572 56500
rect 138 56380 1572 56414
rect 138 56294 1572 56328
rect 138 56208 1572 56242
rect 138 56122 1572 56156
rect 138 56036 1572 56070
rect 138 55950 1572 55984
rect 138 55864 1572 55898
rect 138 55778 1572 55812
rect 138 55692 1572 55726
rect 138 55606 1572 55640
rect 138 55520 1572 55554
rect 138 55434 1572 55468
rect 138 55348 1572 55382
rect 138 55262 1572 55296
rect 138 55176 1572 55210
rect 138 55090 1572 55124
rect 138 55004 1572 55038
rect 138 54918 1572 54952
rect 138 54832 1572 54866
rect 138 54746 1572 54780
rect 138 54660 1572 54694
rect 138 54574 1572 54608
rect 138 54488 1572 54522
rect 138 54402 1572 54436
rect 138 54316 1572 54350
rect 138 54230 1572 54264
rect 138 54144 1572 54178
rect 138 54058 1572 54092
rect 138 53972 1572 54006
rect 138 53886 1572 53920
rect 138 53800 1572 53834
rect 138 53714 1572 53748
rect 138 53628 1572 53662
rect 138 53542 1572 53576
rect 138 53456 1572 53490
rect 138 53370 1572 53404
rect 138 53284 1572 53318
rect 138 53198 1572 53232
rect 138 53112 1572 53146
rect 138 53026 1572 53060
rect 138 52940 1572 52974
rect 138 52854 1572 52888
rect 138 52768 1572 52802
rect 138 52682 1572 52716
rect 138 52596 1572 52630
rect 138 52510 1572 52544
rect 138 52424 1572 52458
rect 138 52338 1572 52372
rect 138 52252 1572 52286
rect 138 52166 1572 52200
rect 138 52080 1572 52114
rect 138 51994 1572 52028
rect 138 51908 1572 51942
rect 138 51822 1572 51856
rect 138 51736 1572 51770
rect 138 51650 1572 51684
rect 138 51564 1572 51598
rect 138 51478 1572 51512
rect 138 51392 1572 51426
rect 138 51306 1572 51340
rect 138 51220 1572 51254
rect 138 51134 1572 51168
rect 138 51048 1572 51082
rect 138 50962 1572 50996
rect 138 50876 1572 50910
rect 138 50790 1572 50824
rect 138 50704 1572 50738
rect 138 50618 1572 50652
rect 138 50532 1572 50566
rect 138 50446 1572 50480
rect 138 50360 1572 50394
rect 138 50274 1572 50308
rect 138 50188 1572 50222
rect 138 50102 1572 50136
rect 138 50016 1572 50050
rect 138 49930 1572 49964
rect 138 49844 1572 49878
rect 138 49758 1572 49792
rect 138 49672 1572 49706
rect 138 49586 1572 49620
rect 138 49500 1572 49534
rect 138 49414 1572 49448
rect 138 49328 1572 49362
rect 138 49242 1572 49276
rect 138 49156 1572 49190
rect 138 49070 1572 49104
rect 138 48984 1572 49018
rect 138 48898 1572 48932
rect 138 48812 1572 48846
rect 138 48726 1572 48760
rect 138 48640 1572 48674
rect 138 48554 1572 48588
rect 138 48468 1572 48502
rect 138 48382 1572 48416
rect 138 48296 1572 48330
rect 138 48210 1572 48244
rect 138 48124 1572 48158
rect 138 48038 1572 48072
rect 138 47952 1572 47986
rect 138 47866 1572 47900
rect 138 47780 1572 47814
rect 138 47694 1572 47728
rect 138 47608 1572 47642
rect 138 47522 1572 47556
rect 138 47436 1572 47470
rect 138 47350 1572 47384
rect 138 47264 1572 47298
rect 138 47178 1572 47212
rect 138 47092 1572 47126
rect 138 47006 1572 47040
rect 138 46920 1572 46954
rect 138 46834 1572 46868
rect 138 46748 1572 46782
rect 138 46662 1572 46696
rect 138 46576 1572 46610
rect 138 46490 1572 46524
rect 138 46404 1572 46438
rect 138 46318 1572 46352
rect 138 46232 1572 46266
rect 138 46146 1572 46180
rect 138 46060 1572 46094
rect 138 45974 1572 46008
rect 138 45888 1572 45922
rect 138 45802 1572 45836
rect 138 45716 1572 45750
rect 138 45630 1572 45664
rect 138 45544 1572 45578
rect 138 45458 1572 45492
rect 138 45372 1572 45406
rect 138 45286 1572 45320
rect 138 45200 1572 45234
rect 138 45114 1572 45148
rect 138 45028 1572 45062
rect 138 44942 1572 44976
rect 138 44856 1572 44890
rect 138 44770 1572 44804
rect 138 44684 1572 44718
rect 138 44598 1572 44632
rect 138 44512 1572 44546
rect 138 44426 1572 44460
rect 138 44340 1572 44374
rect 138 44254 1572 44288
rect 138 44168 1572 44202
rect 138 44082 1572 44116
rect 138 43996 1572 44030
rect 138 43910 1572 43944
rect 138 43824 1572 43858
rect 138 43738 1572 43772
rect 138 43652 1572 43686
rect 138 43566 1572 43600
rect 138 43480 1572 43514
rect 138 43394 1572 43428
rect 138 43308 1572 43342
rect 138 43222 1572 43256
rect 138 43136 1572 43170
rect 138 43050 1572 43084
rect 138 42964 1572 42998
rect 138 42878 1572 42912
rect 138 42792 1572 42826
rect 138 42706 1572 42740
rect 138 42620 1572 42654
rect 138 42534 1572 42568
rect 138 42448 1572 42482
rect 138 42362 1572 42396
rect 138 42276 1572 42310
rect 138 42190 1572 42224
rect 138 42104 1572 42138
rect 138 42018 1572 42052
rect 138 41932 1572 41966
rect 138 41846 1572 41880
rect 138 41760 1572 41794
rect 138 41674 1572 41708
rect 138 41588 1572 41622
rect 138 41502 1572 41536
rect 138 41416 1572 41450
rect 138 41330 1572 41364
rect 138 41244 1572 41278
rect 138 41158 1572 41192
rect 138 41072 1572 41106
rect 138 40986 1572 41020
rect 138 40900 1572 40934
rect 138 40814 1572 40848
rect 138 40728 1572 40762
rect 138 40642 1572 40676
rect 138 40556 1572 40590
rect 138 40470 1572 40504
rect 138 40384 1572 40418
rect 138 40298 1572 40332
rect 138 40212 1572 40246
rect 138 40126 1572 40160
rect 138 40040 1572 40074
rect 138 39954 1572 39988
rect 138 39868 1572 39902
rect 138 39782 1572 39816
rect 138 39696 1572 39730
rect 138 39610 1572 39644
rect 138 39524 1572 39558
rect 138 39438 1572 39472
rect 138 39352 1572 39386
rect 138 39266 1572 39300
rect 138 39180 1572 39214
rect 138 39094 1572 39128
rect 138 39008 1572 39042
rect 138 38922 1572 38956
rect 138 38836 1572 38870
rect 138 38750 1572 38784
rect 138 38664 1572 38698
rect 138 38578 1572 38612
rect 138 38492 1572 38526
rect 138 38406 1572 38440
rect 138 38320 1572 38354
rect 138 38234 1572 38268
rect 138 38148 1572 38182
rect 138 38062 1572 38096
rect 138 37976 1572 38010
rect 138 37890 1572 37924
rect 138 37804 1572 37838
rect 138 37718 1572 37752
rect 138 37632 1572 37666
rect 138 37546 1572 37580
rect 138 37460 1572 37494
rect 138 37374 1572 37408
rect 138 37288 1572 37322
rect 138 37202 1572 37236
rect 138 37116 1572 37150
rect 138 37030 1572 37064
rect 138 36944 1572 36978
rect 138 36858 1572 36892
rect 138 36772 1572 36806
rect 138 36686 1572 36720
rect 138 36600 1572 36634
rect 138 36514 1572 36548
rect 138 36428 1572 36462
rect 138 36342 1572 36376
rect 138 36256 1572 36290
rect 138 36170 1572 36204
rect 138 36084 1572 36118
rect 138 35998 1572 36032
rect 138 35912 1572 35946
rect 138 35826 1572 35860
rect 138 35740 1572 35774
rect 138 35654 1572 35688
rect 138 35568 1572 35602
rect 138 35482 1572 35516
rect 138 35396 1572 35430
rect 138 35310 1572 35344
rect 138 35224 1572 35258
rect 138 35138 1572 35172
rect 138 35052 1572 35086
rect 138 34966 1572 35000
rect 138 34880 1572 34914
rect 138 34794 1572 34828
rect 138 34708 1572 34742
rect 138 34622 1572 34656
rect 138 34536 1572 34570
rect 138 34450 1572 34484
rect 138 34364 1572 34398
rect 138 34278 1572 34312
rect 138 34192 1572 34226
rect 138 34106 1572 34140
rect 138 34020 1572 34054
rect 138 33934 1572 33968
rect 138 33848 1572 33882
rect 138 33762 1572 33796
rect 138 33676 1572 33710
rect 138 33590 1572 33624
rect 138 33504 1572 33538
rect 138 33418 1572 33452
rect 138 33332 1572 33366
rect 138 33246 1572 33280
rect 138 33160 1572 33194
rect 138 33074 1572 33108
rect 138 32988 1572 33022
rect 138 32902 1572 32936
rect 138 32816 1572 32850
rect 138 32730 1572 32764
rect 138 32644 1572 32678
rect 138 32558 1572 32592
rect 138 32472 1572 32506
rect 138 32386 1572 32420
rect 138 32300 1572 32334
rect 138 32214 1572 32248
rect 138 32128 1572 32162
rect 138 32042 1572 32076
rect 138 31956 1572 31990
rect 138 31870 1572 31904
rect 138 31784 1572 31818
rect 138 31698 1572 31732
rect 138 31612 1572 31646
rect 138 31526 1572 31560
rect 138 31440 1572 31474
rect 138 31354 1572 31388
rect 138 31268 1572 31302
rect 138 31182 1572 31216
rect 138 31096 1572 31130
rect 138 31010 1572 31044
rect 138 30924 1572 30958
rect 138 30838 1572 30872
rect 138 30752 1572 30786
rect 138 30666 1572 30700
rect 138 30580 1572 30614
rect 138 30494 1572 30528
rect 138 30408 1572 30442
rect 138 30322 1572 30356
rect 138 30236 1572 30270
rect 138 30150 1572 30184
rect 138 30064 1572 30098
rect 138 29978 1572 30012
rect 138 29892 1572 29926
rect 138 29806 1572 29840
rect 138 29720 1572 29754
rect 138 29634 1572 29668
rect 138 29548 1572 29582
rect 138 29462 1572 29496
rect 138 29376 1572 29410
rect 138 29290 1572 29324
rect 138 29204 1572 29238
rect 138 29118 1572 29152
rect 138 29032 1572 29066
rect 138 28946 1572 28980
rect 138 28860 1572 28894
rect 138 28774 1572 28808
rect 138 28688 1572 28722
rect 138 28602 1572 28636
rect 138 28516 1572 28550
rect 138 28430 1572 28464
rect 138 28344 1572 28378
rect 138 28258 1572 28292
rect 138 28172 1572 28206
rect 138 28086 1572 28120
rect 138 28000 1572 28034
rect 138 27914 1572 27948
rect 138 27828 1572 27862
rect 138 27742 1572 27776
rect 138 27656 1572 27690
rect 138 27570 1572 27604
rect 138 27484 1572 27518
rect 138 27398 1572 27432
rect 138 27312 1572 27346
rect 138 27226 1572 27260
rect 138 27140 1572 27174
rect 138 27054 1572 27088
rect 138 26968 1572 27002
rect 138 26882 1572 26916
rect 138 26796 1572 26830
rect 138 26710 1572 26744
rect 138 26624 1572 26658
rect 138 26538 1572 26572
rect 138 26452 1572 26486
rect 138 26366 1572 26400
rect 138 26280 1572 26314
rect 138 26194 1572 26228
rect 138 26108 1572 26142
rect 138 26022 1572 26056
rect 138 25936 1572 25970
rect 138 25850 1572 25884
rect 138 25764 1572 25798
rect 138 25678 1572 25712
rect 138 25592 1572 25626
rect 138 25506 1572 25540
rect 138 25420 1572 25454
rect 138 25334 1572 25368
rect 138 25248 1572 25282
rect 138 25162 1572 25196
rect 138 25076 1572 25110
rect 138 24990 1572 25024
rect 138 24904 1572 24938
rect 138 24818 1572 24852
rect 138 24732 1572 24766
rect 138 24646 1572 24680
rect 138 24560 1572 24594
rect 138 24474 1572 24508
rect 138 24388 1572 24422
rect 138 24302 1572 24336
rect 138 24216 1572 24250
rect 138 24130 1572 24164
rect 138 24044 1572 24078
rect 138 23958 1572 23992
rect 138 23872 1572 23906
rect 138 23786 1572 23820
rect 138 23700 1572 23734
rect 138 23614 1572 23648
rect 138 23528 1572 23562
rect 138 23442 1572 23476
rect 138 23356 1572 23390
rect 138 23270 1572 23304
rect 138 23184 1572 23218
rect 138 23098 1572 23132
rect 138 23012 1572 23046
rect 138 22926 1572 22960
rect 138 22840 1572 22874
rect 138 22754 1572 22788
rect 138 22668 1572 22702
rect 138 22582 1572 22616
rect 138 22496 1572 22530
rect 138 22410 1572 22444
rect 138 22324 1572 22358
rect 138 22238 1572 22272
rect 138 22152 1572 22186
rect 138 22066 1572 22100
rect 138 21980 1572 22014
rect 138 21894 1572 21928
rect 138 21808 1572 21842
rect 138 21722 1572 21756
rect 138 21636 1572 21670
rect 138 21550 1572 21584
rect 138 21464 1572 21498
rect 138 21378 1572 21412
rect 138 21292 1572 21326
rect 138 21206 1572 21240
rect 138 21120 1572 21154
rect 138 21034 1572 21068
rect 138 20948 1572 20982
rect 138 20862 1572 20896
rect 138 20776 1572 20810
rect 138 20690 1572 20724
rect 138 20604 1572 20638
rect 138 20518 1572 20552
rect 138 20432 1572 20466
rect 138 20346 1572 20380
rect 138 20260 1572 20294
rect 138 20174 1572 20208
rect 138 20088 1572 20122
rect 138 20002 1572 20036
rect 138 19916 1572 19950
rect 138 19830 1572 19864
rect 138 19744 1572 19778
rect 138 19658 1572 19692
rect 138 19572 1572 19606
rect 138 19486 1572 19520
rect 138 19400 1572 19434
rect 138 19314 1572 19348
rect 138 19228 1572 19262
rect 138 19142 1572 19176
rect 138 19056 1572 19090
rect 138 18970 1572 19004
rect 138 18884 1572 18918
rect 138 18798 1572 18832
rect 138 18712 1572 18746
rect 138 18626 1572 18660
rect 138 18540 1572 18574
rect 138 18454 1572 18488
rect 138 18368 1572 18402
rect 138 18282 1572 18316
rect 138 18196 1572 18230
rect 138 18110 1572 18144
rect 138 18024 1572 18058
rect 138 17938 1572 17972
rect 138 17852 1572 17886
rect 138 17766 1572 17800
rect 138 17680 1572 17714
rect 138 17594 1572 17628
rect 138 17508 1572 17542
rect 138 17422 1572 17456
rect 138 17336 1572 17370
rect 138 17250 1572 17284
rect 138 17164 1572 17198
rect 138 17078 1572 17112
rect 138 16992 1572 17026
rect 138 16906 1572 16940
rect 138 16820 1572 16854
rect 138 16734 1572 16768
rect 138 16648 1572 16682
rect 138 16562 1572 16596
rect 138 16476 1572 16510
rect 138 16390 1572 16424
rect 138 16304 1572 16338
rect 138 16218 1572 16252
rect 138 16132 1572 16166
rect 138 16046 1572 16080
rect 138 15960 1572 15994
rect 138 15874 1572 15908
rect 138 15788 1572 15822
rect 138 15702 1572 15736
rect 138 15616 1572 15650
rect 138 15530 1572 15564
rect 138 15444 1572 15478
rect 138 15358 1572 15392
rect 138 15272 1572 15306
rect 138 15186 1572 15220
rect 138 15100 1572 15134
rect 138 15014 1572 15048
rect 138 14928 1572 14962
rect 138 14842 1572 14876
rect 138 14756 1572 14790
rect 138 14670 1572 14704
rect 138 14584 1572 14618
rect 138 14498 1572 14532
rect 138 14412 1572 14446
rect 138 14326 1572 14360
rect 138 14240 1572 14274
rect 138 14154 1572 14188
rect 138 14068 1572 14102
rect 138 13982 1572 14016
rect 138 13896 1572 13930
rect 138 13810 1572 13844
rect 138 13724 1572 13758
rect 138 13638 1572 13672
rect 138 13552 1572 13586
rect 138 13466 1572 13500
rect 138 13380 1572 13414
rect 138 13294 1572 13328
rect 138 13208 1572 13242
rect 138 13122 1572 13156
rect 138 13036 1572 13070
rect 138 12950 1572 12984
rect 138 12864 1572 12898
rect 138 12778 1572 12812
rect 138 12692 1572 12726
rect 138 12606 1572 12640
rect 138 12520 1572 12554
rect 138 12434 1572 12468
rect 138 12348 1572 12382
rect 138 12262 1572 12296
rect 138 12176 1572 12210
rect 138 12090 1572 12124
rect 138 12004 1572 12038
rect 138 11918 1572 11952
rect 138 11832 1572 11866
rect 138 11746 1572 11780
rect 138 11660 1572 11694
rect 138 11574 1572 11608
rect 138 11488 1572 11522
rect 138 11402 1572 11436
rect 138 11316 1572 11350
rect 138 11230 1572 11264
rect 138 11144 1572 11178
rect 138 11058 1572 11092
rect 138 10972 1572 11006
rect 138 10886 1572 10920
rect 138 10800 1572 10834
rect 138 10714 1572 10748
rect 138 10628 1572 10662
rect 138 10542 1572 10576
rect 138 10456 1572 10490
rect 138 10370 1572 10404
rect 138 10284 1572 10318
rect 138 10198 1572 10232
rect 138 10112 1572 10146
rect 138 10026 1572 10060
rect 138 9940 1572 9974
rect 138 9854 1572 9888
rect 138 9768 1572 9802
rect 138 9682 1572 9716
rect 138 9596 1572 9630
rect 138 9510 1572 9544
rect 138 9424 1572 9458
rect 138 9338 1572 9372
rect 138 9252 1572 9286
rect 138 9166 1572 9200
rect 138 9080 1572 9114
rect 138 8994 1572 9028
rect 138 8908 1572 8942
rect 138 8822 1572 8856
rect 138 8736 1572 8770
rect 138 8650 1572 8684
rect 138 8564 1572 8598
rect 138 8478 1572 8512
rect 138 8392 1572 8426
rect 138 8306 1572 8340
rect 138 8220 1572 8254
rect 138 8134 1572 8168
rect 138 8048 1572 8082
rect 138 7962 1572 7996
rect 138 7876 1572 7910
rect 138 7790 1572 7824
rect 138 7704 1572 7738
rect 138 7618 1572 7652
rect 138 7532 1572 7566
rect 138 7446 1572 7480
rect 138 7360 1572 7394
rect 138 7274 1572 7308
rect 138 7188 1572 7222
rect 138 7102 1572 7136
rect 138 7016 1572 7050
rect 138 6930 1572 6964
rect 138 6844 1572 6878
rect 138 6758 1572 6792
rect 138 6672 1572 6706
rect 138 6586 1572 6620
rect 138 6500 1572 6534
rect 138 6414 1572 6448
rect 138 6328 1572 6362
rect 138 6242 1572 6276
rect 138 6156 1572 6190
rect 138 6070 1572 6104
rect 138 5984 1572 6018
rect 138 5898 1572 5932
rect 138 5812 1572 5846
rect 138 5726 1572 5760
rect 138 5640 1572 5674
rect 138 5554 1572 5588
rect 138 5468 1572 5502
rect 138 5382 1572 5416
rect 138 5296 1572 5330
rect 138 5210 1572 5244
rect 138 5124 1572 5158
rect 138 5038 1572 5072
rect 138 4952 1572 4986
rect 138 4866 1572 4900
rect 138 4780 1572 4814
rect 138 4694 1572 4728
rect 138 4608 1572 4642
rect 138 4522 1572 4556
rect 138 4436 1572 4470
rect 138 4350 1572 4384
rect 138 4264 1572 4298
rect 138 4178 1572 4212
rect 138 4092 1572 4126
rect 138 4006 1572 4040
rect 138 3920 1572 3954
rect 138 3834 1572 3868
rect 138 3748 1572 3782
rect 138 3662 1572 3696
rect 138 3576 1572 3610
rect 138 3490 1572 3524
rect 138 3404 1572 3438
rect 138 3318 1572 3352
rect 138 3232 1572 3266
rect 138 3146 1572 3180
rect 138 3060 1572 3094
rect 138 2974 1572 3008
rect 138 2888 1572 2922
rect 138 2802 1572 2836
rect 138 2716 1572 2750
rect 138 2630 1572 2664
rect 138 2544 1572 2578
rect 138 2458 1572 2492
rect 138 2372 1572 2406
rect 138 2286 1572 2320
rect 138 2200 1572 2234
rect 138 2114 1572 2148
rect 138 2028 1572 2062
rect 138 1942 1572 1976
rect 138 1856 1572 1890
rect 138 1770 1572 1804
rect 138 1684 1572 1718
rect 138 1598 1572 1632
rect 138 1512 1572 1546
rect 138 1426 1572 1460
rect 138 1340 1572 1374
rect 138 1254 1572 1288
rect 138 1168 1572 1202
rect 138 1082 1572 1116
rect 138 996 1572 1030
rect 138 910 1572 944
rect 138 824 1572 858
rect 138 738 1572 772
rect 138 652 1572 686
rect 138 566 1572 600
rect 138 480 1572 514
rect 138 394 1572 428
rect 138 308 1572 342
rect 138 222 1572 256
rect 138 136 1572 170
<< nsubdiff >>
rect 36 100168 100 100202
rect 1680 100168 1744 100202
rect 36 100138 70 100168
rect 1710 100138 1744 100168
rect 36 70 70 100
rect 1710 70 1744 100
rect 36 36 100 70
rect 1680 36 1744 70
<< nsubdiffcont >>
rect 100 100168 1680 100202
rect 36 100 70 100138
rect 1710 100 1744 100138
rect 100 36 1680 70
<< poly >>
rect 1618 100059 1672 100075
rect 1618 100057 1628 100059
rect 104 100027 130 100057
rect 1580 100027 1628 100057
rect 1618 99971 1628 100027
rect 104 99941 130 99971
rect 1580 99941 1628 99971
rect 1618 99885 1628 99941
rect 104 99855 130 99885
rect 1580 99855 1628 99885
rect 1618 99799 1628 99855
rect 104 99769 130 99799
rect 1580 99769 1628 99799
rect 1618 99713 1628 99769
rect 104 99683 130 99713
rect 1580 99683 1628 99713
rect 1618 99627 1628 99683
rect 104 99597 130 99627
rect 1580 99597 1628 99627
rect 1618 99541 1628 99597
rect 104 99511 130 99541
rect 1580 99511 1628 99541
rect 1618 99455 1628 99511
rect 104 99425 130 99455
rect 1580 99425 1628 99455
rect 1618 99369 1628 99425
rect 104 99339 130 99369
rect 1580 99339 1628 99369
rect 1618 99283 1628 99339
rect 104 99253 130 99283
rect 1580 99253 1628 99283
rect 1618 99197 1628 99253
rect 104 99167 130 99197
rect 1580 99167 1628 99197
rect 1618 99111 1628 99167
rect 104 99081 130 99111
rect 1580 99081 1628 99111
rect 1618 99025 1628 99081
rect 104 98995 130 99025
rect 1580 98995 1628 99025
rect 1618 98939 1628 98995
rect 104 98909 130 98939
rect 1580 98909 1628 98939
rect 1618 98853 1628 98909
rect 104 98823 130 98853
rect 1580 98823 1628 98853
rect 1618 98767 1628 98823
rect 104 98737 130 98767
rect 1580 98737 1628 98767
rect 1618 98681 1628 98737
rect 104 98651 130 98681
rect 1580 98651 1628 98681
rect 1618 98595 1628 98651
rect 104 98565 130 98595
rect 1580 98565 1628 98595
rect 1618 98509 1628 98565
rect 104 98479 130 98509
rect 1580 98479 1628 98509
rect 1618 98423 1628 98479
rect 104 98393 130 98423
rect 1580 98393 1628 98423
rect 1618 98337 1628 98393
rect 104 98307 130 98337
rect 1580 98307 1628 98337
rect 1618 98251 1628 98307
rect 104 98221 130 98251
rect 1580 98221 1628 98251
rect 1618 98165 1628 98221
rect 104 98135 130 98165
rect 1580 98135 1628 98165
rect 1618 98079 1628 98135
rect 104 98049 130 98079
rect 1580 98049 1628 98079
rect 1618 97993 1628 98049
rect 104 97963 130 97993
rect 1580 97963 1628 97993
rect 1618 97907 1628 97963
rect 104 97877 130 97907
rect 1580 97877 1628 97907
rect 1618 97821 1628 97877
rect 104 97791 130 97821
rect 1580 97791 1628 97821
rect 1618 97735 1628 97791
rect 104 97705 130 97735
rect 1580 97705 1628 97735
rect 1618 97649 1628 97705
rect 104 97619 130 97649
rect 1580 97619 1628 97649
rect 1618 97563 1628 97619
rect 104 97533 130 97563
rect 1580 97533 1628 97563
rect 1618 97477 1628 97533
rect 104 97447 130 97477
rect 1580 97447 1628 97477
rect 1618 97391 1628 97447
rect 104 97361 130 97391
rect 1580 97361 1628 97391
rect 1618 97305 1628 97361
rect 104 97275 130 97305
rect 1580 97275 1628 97305
rect 1618 97219 1628 97275
rect 104 97189 130 97219
rect 1580 97189 1628 97219
rect 1618 97133 1628 97189
rect 104 97103 130 97133
rect 1580 97103 1628 97133
rect 1618 97047 1628 97103
rect 104 97017 130 97047
rect 1580 97017 1628 97047
rect 1618 96961 1628 97017
rect 104 96931 130 96961
rect 1580 96931 1628 96961
rect 1618 96875 1628 96931
rect 104 96845 130 96875
rect 1580 96845 1628 96875
rect 1618 96789 1628 96845
rect 104 96759 130 96789
rect 1580 96759 1628 96789
rect 1618 96703 1628 96759
rect 104 96673 130 96703
rect 1580 96673 1628 96703
rect 1618 96617 1628 96673
rect 104 96587 130 96617
rect 1580 96587 1628 96617
rect 1618 96531 1628 96587
rect 104 96501 130 96531
rect 1580 96501 1628 96531
rect 1618 96445 1628 96501
rect 104 96415 130 96445
rect 1580 96415 1628 96445
rect 1618 96359 1628 96415
rect 104 96329 130 96359
rect 1580 96329 1628 96359
rect 1618 96273 1628 96329
rect 104 96243 130 96273
rect 1580 96243 1628 96273
rect 1618 96187 1628 96243
rect 104 96157 130 96187
rect 1580 96157 1628 96187
rect 1618 96101 1628 96157
rect 104 96071 130 96101
rect 1580 96071 1628 96101
rect 1618 96015 1628 96071
rect 104 95985 130 96015
rect 1580 95985 1628 96015
rect 1618 95929 1628 95985
rect 104 95899 130 95929
rect 1580 95899 1628 95929
rect 1618 95843 1628 95899
rect 104 95813 130 95843
rect 1580 95813 1628 95843
rect 1618 95757 1628 95813
rect 104 95727 130 95757
rect 1580 95727 1628 95757
rect 1618 95671 1628 95727
rect 104 95641 130 95671
rect 1580 95641 1628 95671
rect 1618 95585 1628 95641
rect 104 95555 130 95585
rect 1580 95555 1628 95585
rect 1618 95499 1628 95555
rect 104 95469 130 95499
rect 1580 95469 1628 95499
rect 1618 95413 1628 95469
rect 104 95383 130 95413
rect 1580 95383 1628 95413
rect 1618 95327 1628 95383
rect 104 95297 130 95327
rect 1580 95297 1628 95327
rect 1618 95241 1628 95297
rect 104 95211 130 95241
rect 1580 95211 1628 95241
rect 1618 95155 1628 95211
rect 104 95125 130 95155
rect 1580 95125 1628 95155
rect 1618 95069 1628 95125
rect 104 95039 130 95069
rect 1580 95039 1628 95069
rect 1618 94983 1628 95039
rect 104 94953 130 94983
rect 1580 94953 1628 94983
rect 1618 94897 1628 94953
rect 104 94867 130 94897
rect 1580 94867 1628 94897
rect 1618 94811 1628 94867
rect 104 94781 130 94811
rect 1580 94781 1628 94811
rect 1618 94725 1628 94781
rect 104 94695 130 94725
rect 1580 94695 1628 94725
rect 1618 94639 1628 94695
rect 104 94609 130 94639
rect 1580 94609 1628 94639
rect 1618 94553 1628 94609
rect 104 94523 130 94553
rect 1580 94523 1628 94553
rect 1618 94467 1628 94523
rect 104 94437 130 94467
rect 1580 94437 1628 94467
rect 1618 94381 1628 94437
rect 104 94351 130 94381
rect 1580 94351 1628 94381
rect 1618 94295 1628 94351
rect 104 94265 130 94295
rect 1580 94265 1628 94295
rect 1618 94209 1628 94265
rect 104 94179 130 94209
rect 1580 94179 1628 94209
rect 1618 94123 1628 94179
rect 104 94093 130 94123
rect 1580 94093 1628 94123
rect 1618 94037 1628 94093
rect 104 94007 130 94037
rect 1580 94007 1628 94037
rect 1618 93951 1628 94007
rect 104 93921 130 93951
rect 1580 93921 1628 93951
rect 1618 93865 1628 93921
rect 104 93835 130 93865
rect 1580 93835 1628 93865
rect 1618 93779 1628 93835
rect 104 93749 130 93779
rect 1580 93749 1628 93779
rect 1618 93693 1628 93749
rect 104 93663 130 93693
rect 1580 93663 1628 93693
rect 1618 93607 1628 93663
rect 104 93577 130 93607
rect 1580 93577 1628 93607
rect 1618 93521 1628 93577
rect 104 93491 130 93521
rect 1580 93491 1628 93521
rect 1618 93435 1628 93491
rect 104 93405 130 93435
rect 1580 93405 1628 93435
rect 1618 93349 1628 93405
rect 104 93319 130 93349
rect 1580 93319 1628 93349
rect 1618 93263 1628 93319
rect 104 93233 130 93263
rect 1580 93233 1628 93263
rect 1618 93177 1628 93233
rect 104 93147 130 93177
rect 1580 93147 1628 93177
rect 1618 93091 1628 93147
rect 104 93061 130 93091
rect 1580 93061 1628 93091
rect 1618 93005 1628 93061
rect 104 92975 130 93005
rect 1580 92975 1628 93005
rect 1618 92919 1628 92975
rect 104 92889 130 92919
rect 1580 92889 1628 92919
rect 1618 92833 1628 92889
rect 104 92803 130 92833
rect 1580 92803 1628 92833
rect 1618 92747 1628 92803
rect 104 92717 130 92747
rect 1580 92717 1628 92747
rect 1618 92661 1628 92717
rect 104 92631 130 92661
rect 1580 92631 1628 92661
rect 1618 92575 1628 92631
rect 104 92545 130 92575
rect 1580 92545 1628 92575
rect 1618 92489 1628 92545
rect 104 92459 130 92489
rect 1580 92459 1628 92489
rect 1618 92403 1628 92459
rect 104 92373 130 92403
rect 1580 92373 1628 92403
rect 1618 92317 1628 92373
rect 104 92287 130 92317
rect 1580 92287 1628 92317
rect 1618 92231 1628 92287
rect 104 92201 130 92231
rect 1580 92201 1628 92231
rect 1618 92145 1628 92201
rect 104 92115 130 92145
rect 1580 92115 1628 92145
rect 1618 92059 1628 92115
rect 104 92029 130 92059
rect 1580 92029 1628 92059
rect 1618 91973 1628 92029
rect 104 91943 130 91973
rect 1580 91943 1628 91973
rect 1618 91887 1628 91943
rect 104 91857 130 91887
rect 1580 91857 1628 91887
rect 1618 91801 1628 91857
rect 104 91771 130 91801
rect 1580 91771 1628 91801
rect 1618 91715 1628 91771
rect 104 91685 130 91715
rect 1580 91685 1628 91715
rect 1618 91629 1628 91685
rect 104 91599 130 91629
rect 1580 91599 1628 91629
rect 1618 91543 1628 91599
rect 104 91513 130 91543
rect 1580 91513 1628 91543
rect 1618 91457 1628 91513
rect 104 91427 130 91457
rect 1580 91427 1628 91457
rect 1618 91371 1628 91427
rect 104 91341 130 91371
rect 1580 91341 1628 91371
rect 1618 91285 1628 91341
rect 104 91255 130 91285
rect 1580 91255 1628 91285
rect 1618 91199 1628 91255
rect 104 91169 130 91199
rect 1580 91169 1628 91199
rect 1618 91113 1628 91169
rect 104 91083 130 91113
rect 1580 91083 1628 91113
rect 1618 91027 1628 91083
rect 104 90997 130 91027
rect 1580 90997 1628 91027
rect 1618 90941 1628 90997
rect 104 90911 130 90941
rect 1580 90911 1628 90941
rect 1618 90855 1628 90911
rect 104 90825 130 90855
rect 1580 90825 1628 90855
rect 1618 90769 1628 90825
rect 104 90739 130 90769
rect 1580 90739 1628 90769
rect 1618 90683 1628 90739
rect 104 90653 130 90683
rect 1580 90653 1628 90683
rect 1618 90597 1628 90653
rect 104 90567 130 90597
rect 1580 90567 1628 90597
rect 1618 90511 1628 90567
rect 104 90481 130 90511
rect 1580 90481 1628 90511
rect 1618 90425 1628 90481
rect 104 90395 130 90425
rect 1580 90395 1628 90425
rect 1618 90339 1628 90395
rect 104 90309 130 90339
rect 1580 90309 1628 90339
rect 1618 90253 1628 90309
rect 104 90223 130 90253
rect 1580 90223 1628 90253
rect 1618 90167 1628 90223
rect 104 90137 130 90167
rect 1580 90137 1628 90167
rect 1618 90081 1628 90137
rect 104 90051 130 90081
rect 1580 90051 1628 90081
rect 1618 89995 1628 90051
rect 104 89965 130 89995
rect 1580 89965 1628 89995
rect 1618 89909 1628 89965
rect 104 89879 130 89909
rect 1580 89879 1628 89909
rect 1618 89823 1628 89879
rect 104 89793 130 89823
rect 1580 89793 1628 89823
rect 1618 89737 1628 89793
rect 104 89707 130 89737
rect 1580 89707 1628 89737
rect 1618 89651 1628 89707
rect 104 89621 130 89651
rect 1580 89621 1628 89651
rect 1618 89565 1628 89621
rect 104 89535 130 89565
rect 1580 89535 1628 89565
rect 1618 89479 1628 89535
rect 104 89449 130 89479
rect 1580 89449 1628 89479
rect 1618 89393 1628 89449
rect 104 89363 130 89393
rect 1580 89363 1628 89393
rect 1618 89307 1628 89363
rect 104 89277 130 89307
rect 1580 89277 1628 89307
rect 1618 89221 1628 89277
rect 104 89191 130 89221
rect 1580 89191 1628 89221
rect 1618 89135 1628 89191
rect 104 89105 130 89135
rect 1580 89105 1628 89135
rect 1618 89049 1628 89105
rect 104 89019 130 89049
rect 1580 89019 1628 89049
rect 1618 88963 1628 89019
rect 104 88933 130 88963
rect 1580 88933 1628 88963
rect 1618 88877 1628 88933
rect 104 88847 130 88877
rect 1580 88847 1628 88877
rect 1618 88791 1628 88847
rect 104 88761 130 88791
rect 1580 88761 1628 88791
rect 1618 88705 1628 88761
rect 104 88675 130 88705
rect 1580 88675 1628 88705
rect 1618 88619 1628 88675
rect 104 88589 130 88619
rect 1580 88589 1628 88619
rect 1618 88533 1628 88589
rect 104 88503 130 88533
rect 1580 88503 1628 88533
rect 1618 88447 1628 88503
rect 104 88417 130 88447
rect 1580 88417 1628 88447
rect 1618 88361 1628 88417
rect 104 88331 130 88361
rect 1580 88331 1628 88361
rect 1618 88275 1628 88331
rect 104 88245 130 88275
rect 1580 88245 1628 88275
rect 1618 88189 1628 88245
rect 104 88159 130 88189
rect 1580 88159 1628 88189
rect 1618 88103 1628 88159
rect 104 88073 130 88103
rect 1580 88073 1628 88103
rect 1618 88017 1628 88073
rect 104 87987 130 88017
rect 1580 87987 1628 88017
rect 1618 87931 1628 87987
rect 104 87901 130 87931
rect 1580 87901 1628 87931
rect 1618 87845 1628 87901
rect 104 87815 130 87845
rect 1580 87815 1628 87845
rect 1618 87759 1628 87815
rect 104 87729 130 87759
rect 1580 87729 1628 87759
rect 1618 87673 1628 87729
rect 104 87643 130 87673
rect 1580 87643 1628 87673
rect 1618 87587 1628 87643
rect 104 87557 130 87587
rect 1580 87557 1628 87587
rect 1618 87501 1628 87557
rect 104 87471 130 87501
rect 1580 87471 1628 87501
rect 1618 87415 1628 87471
rect 104 87385 130 87415
rect 1580 87385 1628 87415
rect 1618 87329 1628 87385
rect 104 87299 130 87329
rect 1580 87299 1628 87329
rect 1618 87243 1628 87299
rect 104 87213 130 87243
rect 1580 87213 1628 87243
rect 1618 87157 1628 87213
rect 104 87127 130 87157
rect 1580 87127 1628 87157
rect 1618 87071 1628 87127
rect 104 87041 130 87071
rect 1580 87041 1628 87071
rect 1618 86985 1628 87041
rect 104 86955 130 86985
rect 1580 86955 1628 86985
rect 1618 86899 1628 86955
rect 104 86869 130 86899
rect 1580 86869 1628 86899
rect 1618 86813 1628 86869
rect 104 86783 130 86813
rect 1580 86783 1628 86813
rect 1618 86727 1628 86783
rect 104 86697 130 86727
rect 1580 86697 1628 86727
rect 1618 86641 1628 86697
rect 104 86611 130 86641
rect 1580 86611 1628 86641
rect 1618 86555 1628 86611
rect 104 86525 130 86555
rect 1580 86525 1628 86555
rect 1618 86469 1628 86525
rect 104 86439 130 86469
rect 1580 86439 1628 86469
rect 1618 86383 1628 86439
rect 104 86353 130 86383
rect 1580 86353 1628 86383
rect 1618 86297 1628 86353
rect 104 86267 130 86297
rect 1580 86267 1628 86297
rect 1618 86211 1628 86267
rect 104 86181 130 86211
rect 1580 86181 1628 86211
rect 1618 86125 1628 86181
rect 104 86095 130 86125
rect 1580 86095 1628 86125
rect 1618 86039 1628 86095
rect 104 86009 130 86039
rect 1580 86009 1628 86039
rect 1618 85953 1628 86009
rect 104 85923 130 85953
rect 1580 85923 1628 85953
rect 1618 85867 1628 85923
rect 104 85837 130 85867
rect 1580 85837 1628 85867
rect 1618 85781 1628 85837
rect 104 85751 130 85781
rect 1580 85751 1628 85781
rect 1618 85695 1628 85751
rect 104 85665 130 85695
rect 1580 85665 1628 85695
rect 1618 85609 1628 85665
rect 104 85579 130 85609
rect 1580 85579 1628 85609
rect 1618 85523 1628 85579
rect 104 85493 130 85523
rect 1580 85493 1628 85523
rect 1618 85437 1628 85493
rect 104 85407 130 85437
rect 1580 85407 1628 85437
rect 1618 85351 1628 85407
rect 104 85321 130 85351
rect 1580 85321 1628 85351
rect 1618 85265 1628 85321
rect 104 85235 130 85265
rect 1580 85235 1628 85265
rect 1618 85179 1628 85235
rect 104 85149 130 85179
rect 1580 85149 1628 85179
rect 1618 85093 1628 85149
rect 104 85063 130 85093
rect 1580 85063 1628 85093
rect 1618 85007 1628 85063
rect 104 84977 130 85007
rect 1580 84977 1628 85007
rect 1618 84921 1628 84977
rect 104 84891 130 84921
rect 1580 84891 1628 84921
rect 1618 84835 1628 84891
rect 104 84805 130 84835
rect 1580 84805 1628 84835
rect 1618 84749 1628 84805
rect 104 84719 130 84749
rect 1580 84719 1628 84749
rect 1618 84663 1628 84719
rect 104 84633 130 84663
rect 1580 84633 1628 84663
rect 1618 84577 1628 84633
rect 104 84547 130 84577
rect 1580 84547 1628 84577
rect 1618 84491 1628 84547
rect 104 84461 130 84491
rect 1580 84461 1628 84491
rect 1618 84405 1628 84461
rect 104 84375 130 84405
rect 1580 84375 1628 84405
rect 1618 84319 1628 84375
rect 104 84289 130 84319
rect 1580 84289 1628 84319
rect 1618 84233 1628 84289
rect 104 84203 130 84233
rect 1580 84203 1628 84233
rect 1618 84147 1628 84203
rect 104 84117 130 84147
rect 1580 84117 1628 84147
rect 1618 84061 1628 84117
rect 104 84031 130 84061
rect 1580 84031 1628 84061
rect 1618 83975 1628 84031
rect 104 83945 130 83975
rect 1580 83945 1628 83975
rect 1618 83889 1628 83945
rect 104 83859 130 83889
rect 1580 83859 1628 83889
rect 1618 83803 1628 83859
rect 104 83773 130 83803
rect 1580 83773 1628 83803
rect 1618 83717 1628 83773
rect 104 83687 130 83717
rect 1580 83687 1628 83717
rect 1618 83631 1628 83687
rect 104 83601 130 83631
rect 1580 83601 1628 83631
rect 1618 83545 1628 83601
rect 104 83515 130 83545
rect 1580 83515 1628 83545
rect 1618 83459 1628 83515
rect 104 83429 130 83459
rect 1580 83429 1628 83459
rect 1618 83373 1628 83429
rect 104 83343 130 83373
rect 1580 83343 1628 83373
rect 1618 83287 1628 83343
rect 104 83257 130 83287
rect 1580 83257 1628 83287
rect 1618 83201 1628 83257
rect 104 83171 130 83201
rect 1580 83171 1628 83201
rect 1618 83115 1628 83171
rect 104 83085 130 83115
rect 1580 83085 1628 83115
rect 1618 83029 1628 83085
rect 104 82999 130 83029
rect 1580 82999 1628 83029
rect 1618 82943 1628 82999
rect 104 82913 130 82943
rect 1580 82913 1628 82943
rect 1618 82857 1628 82913
rect 104 82827 130 82857
rect 1580 82827 1628 82857
rect 1618 82771 1628 82827
rect 104 82741 130 82771
rect 1580 82741 1628 82771
rect 1618 82685 1628 82741
rect 104 82655 130 82685
rect 1580 82655 1628 82685
rect 1618 82599 1628 82655
rect 104 82569 130 82599
rect 1580 82569 1628 82599
rect 1618 82513 1628 82569
rect 104 82483 130 82513
rect 1580 82483 1628 82513
rect 1618 82427 1628 82483
rect 104 82397 130 82427
rect 1580 82397 1628 82427
rect 1618 82341 1628 82397
rect 104 82311 130 82341
rect 1580 82311 1628 82341
rect 1618 82255 1628 82311
rect 104 82225 130 82255
rect 1580 82225 1628 82255
rect 1618 82169 1628 82225
rect 104 82139 130 82169
rect 1580 82139 1628 82169
rect 1618 82083 1628 82139
rect 104 82053 130 82083
rect 1580 82053 1628 82083
rect 1618 81997 1628 82053
rect 104 81967 130 81997
rect 1580 81967 1628 81997
rect 1618 81911 1628 81967
rect 104 81881 130 81911
rect 1580 81881 1628 81911
rect 1618 81825 1628 81881
rect 104 81795 130 81825
rect 1580 81795 1628 81825
rect 1618 81739 1628 81795
rect 104 81709 130 81739
rect 1580 81709 1628 81739
rect 1618 81653 1628 81709
rect 104 81623 130 81653
rect 1580 81623 1628 81653
rect 1618 81567 1628 81623
rect 104 81537 130 81567
rect 1580 81537 1628 81567
rect 1618 81481 1628 81537
rect 104 81451 130 81481
rect 1580 81451 1628 81481
rect 1618 81395 1628 81451
rect 104 81365 130 81395
rect 1580 81365 1628 81395
rect 1618 81309 1628 81365
rect 104 81279 130 81309
rect 1580 81279 1628 81309
rect 1618 81223 1628 81279
rect 104 81193 130 81223
rect 1580 81193 1628 81223
rect 1618 81137 1628 81193
rect 104 81107 130 81137
rect 1580 81107 1628 81137
rect 1618 81051 1628 81107
rect 104 81021 130 81051
rect 1580 81021 1628 81051
rect 1618 80965 1628 81021
rect 104 80935 130 80965
rect 1580 80935 1628 80965
rect 1618 80879 1628 80935
rect 104 80849 130 80879
rect 1580 80849 1628 80879
rect 1618 80793 1628 80849
rect 104 80763 130 80793
rect 1580 80763 1628 80793
rect 1618 80707 1628 80763
rect 104 80677 130 80707
rect 1580 80677 1628 80707
rect 1618 80621 1628 80677
rect 104 80591 130 80621
rect 1580 80591 1628 80621
rect 1618 80535 1628 80591
rect 104 80505 130 80535
rect 1580 80505 1628 80535
rect 1618 80449 1628 80505
rect 104 80419 130 80449
rect 1580 80419 1628 80449
rect 1618 80363 1628 80419
rect 104 80333 130 80363
rect 1580 80333 1628 80363
rect 1618 80277 1628 80333
rect 104 80247 130 80277
rect 1580 80247 1628 80277
rect 1618 80191 1628 80247
rect 104 80161 130 80191
rect 1580 80161 1628 80191
rect 1618 80105 1628 80161
rect 104 80075 130 80105
rect 1580 80075 1628 80105
rect 1618 80019 1628 80075
rect 104 79989 130 80019
rect 1580 79989 1628 80019
rect 1618 79933 1628 79989
rect 104 79903 130 79933
rect 1580 79903 1628 79933
rect 1618 79847 1628 79903
rect 104 79817 130 79847
rect 1580 79817 1628 79847
rect 1618 79761 1628 79817
rect 104 79731 130 79761
rect 1580 79731 1628 79761
rect 1618 79675 1628 79731
rect 104 79645 130 79675
rect 1580 79645 1628 79675
rect 1618 79589 1628 79645
rect 104 79559 130 79589
rect 1580 79559 1628 79589
rect 1618 79503 1628 79559
rect 104 79473 130 79503
rect 1580 79473 1628 79503
rect 1618 79417 1628 79473
rect 104 79387 130 79417
rect 1580 79387 1628 79417
rect 1618 79331 1628 79387
rect 104 79301 130 79331
rect 1580 79301 1628 79331
rect 1618 79245 1628 79301
rect 104 79215 130 79245
rect 1580 79215 1628 79245
rect 1618 79159 1628 79215
rect 104 79129 130 79159
rect 1580 79129 1628 79159
rect 1618 79073 1628 79129
rect 104 79043 130 79073
rect 1580 79043 1628 79073
rect 1618 78987 1628 79043
rect 104 78957 130 78987
rect 1580 78957 1628 78987
rect 1618 78901 1628 78957
rect 104 78871 130 78901
rect 1580 78871 1628 78901
rect 1618 78815 1628 78871
rect 104 78785 130 78815
rect 1580 78785 1628 78815
rect 1618 78729 1628 78785
rect 104 78699 130 78729
rect 1580 78699 1628 78729
rect 1618 78643 1628 78699
rect 104 78613 130 78643
rect 1580 78613 1628 78643
rect 1618 78557 1628 78613
rect 104 78527 130 78557
rect 1580 78527 1628 78557
rect 1618 78471 1628 78527
rect 104 78441 130 78471
rect 1580 78441 1628 78471
rect 1618 78385 1628 78441
rect 104 78355 130 78385
rect 1580 78355 1628 78385
rect 1618 78299 1628 78355
rect 104 78269 130 78299
rect 1580 78269 1628 78299
rect 1618 78213 1628 78269
rect 104 78183 130 78213
rect 1580 78183 1628 78213
rect 1618 78127 1628 78183
rect 104 78097 130 78127
rect 1580 78097 1628 78127
rect 1618 78041 1628 78097
rect 104 78011 130 78041
rect 1580 78011 1628 78041
rect 1618 77955 1628 78011
rect 104 77925 130 77955
rect 1580 77925 1628 77955
rect 1618 77869 1628 77925
rect 104 77839 130 77869
rect 1580 77839 1628 77869
rect 1618 77783 1628 77839
rect 104 77753 130 77783
rect 1580 77753 1628 77783
rect 1618 77697 1628 77753
rect 104 77667 130 77697
rect 1580 77667 1628 77697
rect 1618 77611 1628 77667
rect 104 77581 130 77611
rect 1580 77581 1628 77611
rect 1618 77525 1628 77581
rect 104 77495 130 77525
rect 1580 77495 1628 77525
rect 1618 77439 1628 77495
rect 104 77409 130 77439
rect 1580 77409 1628 77439
rect 1618 77353 1628 77409
rect 104 77323 130 77353
rect 1580 77323 1628 77353
rect 1618 77267 1628 77323
rect 104 77237 130 77267
rect 1580 77237 1628 77267
rect 1618 77181 1628 77237
rect 104 77151 130 77181
rect 1580 77151 1628 77181
rect 1618 77095 1628 77151
rect 104 77065 130 77095
rect 1580 77065 1628 77095
rect 1618 77009 1628 77065
rect 104 76979 130 77009
rect 1580 76979 1628 77009
rect 1618 76923 1628 76979
rect 104 76893 130 76923
rect 1580 76893 1628 76923
rect 1618 76837 1628 76893
rect 104 76807 130 76837
rect 1580 76807 1628 76837
rect 1618 76751 1628 76807
rect 104 76721 130 76751
rect 1580 76721 1628 76751
rect 1618 76665 1628 76721
rect 104 76635 130 76665
rect 1580 76635 1628 76665
rect 1618 76579 1628 76635
rect 104 76549 130 76579
rect 1580 76549 1628 76579
rect 1618 76493 1628 76549
rect 104 76463 130 76493
rect 1580 76463 1628 76493
rect 1618 76407 1628 76463
rect 104 76377 130 76407
rect 1580 76377 1628 76407
rect 1618 76321 1628 76377
rect 104 76291 130 76321
rect 1580 76291 1628 76321
rect 1618 76235 1628 76291
rect 104 76205 130 76235
rect 1580 76205 1628 76235
rect 1618 76149 1628 76205
rect 104 76119 130 76149
rect 1580 76119 1628 76149
rect 1618 76063 1628 76119
rect 104 76033 130 76063
rect 1580 76033 1628 76063
rect 1618 75977 1628 76033
rect 104 75947 130 75977
rect 1580 75947 1628 75977
rect 1618 75891 1628 75947
rect 104 75861 130 75891
rect 1580 75861 1628 75891
rect 1618 75805 1628 75861
rect 104 75775 130 75805
rect 1580 75775 1628 75805
rect 1618 75719 1628 75775
rect 104 75689 130 75719
rect 1580 75689 1628 75719
rect 1618 75633 1628 75689
rect 104 75603 130 75633
rect 1580 75603 1628 75633
rect 1618 75547 1628 75603
rect 104 75517 130 75547
rect 1580 75517 1628 75547
rect 1618 75461 1628 75517
rect 104 75431 130 75461
rect 1580 75431 1628 75461
rect 1618 75375 1628 75431
rect 104 75345 130 75375
rect 1580 75345 1628 75375
rect 1618 75289 1628 75345
rect 104 75259 130 75289
rect 1580 75259 1628 75289
rect 1618 75203 1628 75259
rect 104 75173 130 75203
rect 1580 75173 1628 75203
rect 1618 75117 1628 75173
rect 104 75087 130 75117
rect 1580 75087 1628 75117
rect 1618 75031 1628 75087
rect 104 75001 130 75031
rect 1580 75001 1628 75031
rect 1618 74945 1628 75001
rect 104 74915 130 74945
rect 1580 74915 1628 74945
rect 1618 74859 1628 74915
rect 104 74829 130 74859
rect 1580 74829 1628 74859
rect 1618 74773 1628 74829
rect 104 74743 130 74773
rect 1580 74743 1628 74773
rect 1618 74687 1628 74743
rect 104 74657 130 74687
rect 1580 74657 1628 74687
rect 1618 74601 1628 74657
rect 104 74571 130 74601
rect 1580 74571 1628 74601
rect 1618 74515 1628 74571
rect 104 74485 130 74515
rect 1580 74485 1628 74515
rect 1618 74429 1628 74485
rect 104 74399 130 74429
rect 1580 74399 1628 74429
rect 1618 74343 1628 74399
rect 104 74313 130 74343
rect 1580 74313 1628 74343
rect 1618 74257 1628 74313
rect 104 74227 130 74257
rect 1580 74227 1628 74257
rect 1618 74171 1628 74227
rect 104 74141 130 74171
rect 1580 74141 1628 74171
rect 1618 74085 1628 74141
rect 104 74055 130 74085
rect 1580 74055 1628 74085
rect 1618 73999 1628 74055
rect 104 73969 130 73999
rect 1580 73969 1628 73999
rect 1618 73913 1628 73969
rect 104 73883 130 73913
rect 1580 73883 1628 73913
rect 1618 73827 1628 73883
rect 104 73797 130 73827
rect 1580 73797 1628 73827
rect 1618 73741 1628 73797
rect 104 73711 130 73741
rect 1580 73711 1628 73741
rect 1618 73655 1628 73711
rect 104 73625 130 73655
rect 1580 73625 1628 73655
rect 1618 73569 1628 73625
rect 104 73539 130 73569
rect 1580 73539 1628 73569
rect 1618 73483 1628 73539
rect 104 73453 130 73483
rect 1580 73453 1628 73483
rect 1618 73397 1628 73453
rect 104 73367 130 73397
rect 1580 73367 1628 73397
rect 1618 73311 1628 73367
rect 104 73281 130 73311
rect 1580 73281 1628 73311
rect 1618 73225 1628 73281
rect 104 73195 130 73225
rect 1580 73195 1628 73225
rect 1618 73139 1628 73195
rect 104 73109 130 73139
rect 1580 73109 1628 73139
rect 1618 73053 1628 73109
rect 104 73023 130 73053
rect 1580 73023 1628 73053
rect 1618 72967 1628 73023
rect 104 72937 130 72967
rect 1580 72937 1628 72967
rect 1618 72881 1628 72937
rect 104 72851 130 72881
rect 1580 72851 1628 72881
rect 1618 72795 1628 72851
rect 104 72765 130 72795
rect 1580 72765 1628 72795
rect 1618 72709 1628 72765
rect 104 72679 130 72709
rect 1580 72679 1628 72709
rect 1618 72623 1628 72679
rect 104 72593 130 72623
rect 1580 72593 1628 72623
rect 1618 72537 1628 72593
rect 104 72507 130 72537
rect 1580 72507 1628 72537
rect 1618 72451 1628 72507
rect 104 72421 130 72451
rect 1580 72421 1628 72451
rect 1618 72365 1628 72421
rect 104 72335 130 72365
rect 1580 72335 1628 72365
rect 1618 72279 1628 72335
rect 104 72249 130 72279
rect 1580 72249 1628 72279
rect 1618 72193 1628 72249
rect 104 72163 130 72193
rect 1580 72163 1628 72193
rect 1618 72107 1628 72163
rect 104 72077 130 72107
rect 1580 72077 1628 72107
rect 1618 72021 1628 72077
rect 104 71991 130 72021
rect 1580 71991 1628 72021
rect 1618 71935 1628 71991
rect 104 71905 130 71935
rect 1580 71905 1628 71935
rect 1618 71849 1628 71905
rect 104 71819 130 71849
rect 1580 71819 1628 71849
rect 1618 71763 1628 71819
rect 104 71733 130 71763
rect 1580 71733 1628 71763
rect 1618 71677 1628 71733
rect 104 71647 130 71677
rect 1580 71647 1628 71677
rect 1618 71591 1628 71647
rect 104 71561 130 71591
rect 1580 71561 1628 71591
rect 1618 71505 1628 71561
rect 104 71475 130 71505
rect 1580 71475 1628 71505
rect 1618 71419 1628 71475
rect 104 71389 130 71419
rect 1580 71389 1628 71419
rect 1618 71333 1628 71389
rect 104 71303 130 71333
rect 1580 71303 1628 71333
rect 1618 71247 1628 71303
rect 104 71217 130 71247
rect 1580 71217 1628 71247
rect 1618 71161 1628 71217
rect 104 71131 130 71161
rect 1580 71131 1628 71161
rect 1618 71075 1628 71131
rect 104 71045 130 71075
rect 1580 71045 1628 71075
rect 1618 70989 1628 71045
rect 104 70959 130 70989
rect 1580 70959 1628 70989
rect 1618 70903 1628 70959
rect 104 70873 130 70903
rect 1580 70873 1628 70903
rect 1618 70817 1628 70873
rect 104 70787 130 70817
rect 1580 70787 1628 70817
rect 1618 70731 1628 70787
rect 104 70701 130 70731
rect 1580 70701 1628 70731
rect 1618 70645 1628 70701
rect 104 70615 130 70645
rect 1580 70615 1628 70645
rect 1618 70559 1628 70615
rect 104 70529 130 70559
rect 1580 70529 1628 70559
rect 1618 70473 1628 70529
rect 104 70443 130 70473
rect 1580 70443 1628 70473
rect 1618 70387 1628 70443
rect 104 70357 130 70387
rect 1580 70357 1628 70387
rect 1618 70301 1628 70357
rect 104 70271 130 70301
rect 1580 70271 1628 70301
rect 1618 70215 1628 70271
rect 104 70185 130 70215
rect 1580 70185 1628 70215
rect 1618 70129 1628 70185
rect 104 70099 130 70129
rect 1580 70099 1628 70129
rect 1618 70043 1628 70099
rect 104 70013 130 70043
rect 1580 70013 1628 70043
rect 1618 69957 1628 70013
rect 104 69927 130 69957
rect 1580 69927 1628 69957
rect 1618 69871 1628 69927
rect 104 69841 130 69871
rect 1580 69841 1628 69871
rect 1618 69785 1628 69841
rect 104 69755 130 69785
rect 1580 69755 1628 69785
rect 1618 69699 1628 69755
rect 104 69669 130 69699
rect 1580 69669 1628 69699
rect 1618 69613 1628 69669
rect 104 69583 130 69613
rect 1580 69583 1628 69613
rect 1618 69527 1628 69583
rect 104 69497 130 69527
rect 1580 69497 1628 69527
rect 1618 69441 1628 69497
rect 104 69411 130 69441
rect 1580 69411 1628 69441
rect 1618 69355 1628 69411
rect 104 69325 130 69355
rect 1580 69325 1628 69355
rect 1618 69269 1628 69325
rect 104 69239 130 69269
rect 1580 69239 1628 69269
rect 1618 69183 1628 69239
rect 104 69153 130 69183
rect 1580 69153 1628 69183
rect 1618 69097 1628 69153
rect 104 69067 130 69097
rect 1580 69067 1628 69097
rect 1618 69011 1628 69067
rect 104 68981 130 69011
rect 1580 68981 1628 69011
rect 1618 68925 1628 68981
rect 104 68895 130 68925
rect 1580 68895 1628 68925
rect 1618 68839 1628 68895
rect 104 68809 130 68839
rect 1580 68809 1628 68839
rect 1618 68753 1628 68809
rect 104 68723 130 68753
rect 1580 68723 1628 68753
rect 1618 68667 1628 68723
rect 104 68637 130 68667
rect 1580 68637 1628 68667
rect 1618 68581 1628 68637
rect 104 68551 130 68581
rect 1580 68551 1628 68581
rect 1618 68495 1628 68551
rect 104 68465 130 68495
rect 1580 68465 1628 68495
rect 1618 68409 1628 68465
rect 104 68379 130 68409
rect 1580 68379 1628 68409
rect 1618 68323 1628 68379
rect 104 68293 130 68323
rect 1580 68293 1628 68323
rect 1618 68237 1628 68293
rect 104 68207 130 68237
rect 1580 68207 1628 68237
rect 1618 68151 1628 68207
rect 104 68121 130 68151
rect 1580 68121 1628 68151
rect 1618 68065 1628 68121
rect 104 68035 130 68065
rect 1580 68035 1628 68065
rect 1618 67979 1628 68035
rect 104 67949 130 67979
rect 1580 67949 1628 67979
rect 1618 67893 1628 67949
rect 104 67863 130 67893
rect 1580 67863 1628 67893
rect 1618 67807 1628 67863
rect 104 67777 130 67807
rect 1580 67777 1628 67807
rect 1618 67721 1628 67777
rect 104 67691 130 67721
rect 1580 67691 1628 67721
rect 1618 67635 1628 67691
rect 104 67605 130 67635
rect 1580 67605 1628 67635
rect 1618 67549 1628 67605
rect 104 67519 130 67549
rect 1580 67519 1628 67549
rect 1618 67463 1628 67519
rect 104 67433 130 67463
rect 1580 67433 1628 67463
rect 1618 67377 1628 67433
rect 104 67347 130 67377
rect 1580 67347 1628 67377
rect 1618 67291 1628 67347
rect 104 67261 130 67291
rect 1580 67261 1628 67291
rect 1618 67205 1628 67261
rect 104 67175 130 67205
rect 1580 67175 1628 67205
rect 1618 67119 1628 67175
rect 104 67089 130 67119
rect 1580 67089 1628 67119
rect 1618 67033 1628 67089
rect 104 67003 130 67033
rect 1580 67003 1628 67033
rect 1618 66947 1628 67003
rect 104 66917 130 66947
rect 1580 66917 1628 66947
rect 1618 66861 1628 66917
rect 104 66831 130 66861
rect 1580 66831 1628 66861
rect 1618 66775 1628 66831
rect 104 66745 130 66775
rect 1580 66745 1628 66775
rect 1618 66689 1628 66745
rect 104 66659 130 66689
rect 1580 66659 1628 66689
rect 1618 66603 1628 66659
rect 104 66573 130 66603
rect 1580 66573 1628 66603
rect 1618 66517 1628 66573
rect 104 66487 130 66517
rect 1580 66487 1628 66517
rect 1618 66431 1628 66487
rect 104 66401 130 66431
rect 1580 66401 1628 66431
rect 1618 66345 1628 66401
rect 104 66315 130 66345
rect 1580 66315 1628 66345
rect 1618 66259 1628 66315
rect 104 66229 130 66259
rect 1580 66229 1628 66259
rect 1618 66173 1628 66229
rect 104 66143 130 66173
rect 1580 66143 1628 66173
rect 1618 66087 1628 66143
rect 104 66057 130 66087
rect 1580 66057 1628 66087
rect 1618 66001 1628 66057
rect 104 65971 130 66001
rect 1580 65971 1628 66001
rect 1618 65915 1628 65971
rect 104 65885 130 65915
rect 1580 65885 1628 65915
rect 1618 65829 1628 65885
rect 104 65799 130 65829
rect 1580 65799 1628 65829
rect 1618 65743 1628 65799
rect 104 65713 130 65743
rect 1580 65713 1628 65743
rect 1618 65657 1628 65713
rect 104 65627 130 65657
rect 1580 65627 1628 65657
rect 1618 65571 1628 65627
rect 104 65541 130 65571
rect 1580 65541 1628 65571
rect 1618 65485 1628 65541
rect 104 65455 130 65485
rect 1580 65455 1628 65485
rect 1618 65399 1628 65455
rect 104 65369 130 65399
rect 1580 65369 1628 65399
rect 1618 65313 1628 65369
rect 104 65283 130 65313
rect 1580 65283 1628 65313
rect 1618 65227 1628 65283
rect 104 65197 130 65227
rect 1580 65197 1628 65227
rect 1618 65141 1628 65197
rect 104 65111 130 65141
rect 1580 65111 1628 65141
rect 1618 65055 1628 65111
rect 104 65025 130 65055
rect 1580 65025 1628 65055
rect 1618 64969 1628 65025
rect 104 64939 130 64969
rect 1580 64939 1628 64969
rect 1618 64883 1628 64939
rect 104 64853 130 64883
rect 1580 64853 1628 64883
rect 1618 64797 1628 64853
rect 104 64767 130 64797
rect 1580 64767 1628 64797
rect 1618 64711 1628 64767
rect 104 64681 130 64711
rect 1580 64681 1628 64711
rect 1618 64625 1628 64681
rect 104 64595 130 64625
rect 1580 64595 1628 64625
rect 1618 64539 1628 64595
rect 104 64509 130 64539
rect 1580 64509 1628 64539
rect 1618 64453 1628 64509
rect 104 64423 130 64453
rect 1580 64423 1628 64453
rect 1618 64367 1628 64423
rect 104 64337 130 64367
rect 1580 64337 1628 64367
rect 1618 64281 1628 64337
rect 104 64251 130 64281
rect 1580 64251 1628 64281
rect 1618 64195 1628 64251
rect 104 64165 130 64195
rect 1580 64165 1628 64195
rect 1618 64109 1628 64165
rect 104 64079 130 64109
rect 1580 64079 1628 64109
rect 1618 64023 1628 64079
rect 104 63993 130 64023
rect 1580 63993 1628 64023
rect 1618 63937 1628 63993
rect 104 63907 130 63937
rect 1580 63907 1628 63937
rect 1618 63851 1628 63907
rect 104 63821 130 63851
rect 1580 63821 1628 63851
rect 1618 63765 1628 63821
rect 104 63735 130 63765
rect 1580 63735 1628 63765
rect 1618 63679 1628 63735
rect 104 63649 130 63679
rect 1580 63649 1628 63679
rect 1618 63593 1628 63649
rect 104 63563 130 63593
rect 1580 63563 1628 63593
rect 1618 63507 1628 63563
rect 104 63477 130 63507
rect 1580 63477 1628 63507
rect 1618 63421 1628 63477
rect 104 63391 130 63421
rect 1580 63391 1628 63421
rect 1618 63335 1628 63391
rect 104 63305 130 63335
rect 1580 63305 1628 63335
rect 1618 63249 1628 63305
rect 104 63219 130 63249
rect 1580 63219 1628 63249
rect 1618 63163 1628 63219
rect 104 63133 130 63163
rect 1580 63133 1628 63163
rect 1618 63077 1628 63133
rect 104 63047 130 63077
rect 1580 63047 1628 63077
rect 1618 62991 1628 63047
rect 104 62961 130 62991
rect 1580 62961 1628 62991
rect 1618 62905 1628 62961
rect 104 62875 130 62905
rect 1580 62875 1628 62905
rect 1618 62819 1628 62875
rect 104 62789 130 62819
rect 1580 62789 1628 62819
rect 1618 62733 1628 62789
rect 104 62703 130 62733
rect 1580 62703 1628 62733
rect 1618 62647 1628 62703
rect 104 62617 130 62647
rect 1580 62617 1628 62647
rect 1618 62561 1628 62617
rect 104 62531 130 62561
rect 1580 62531 1628 62561
rect 1618 62475 1628 62531
rect 104 62445 130 62475
rect 1580 62445 1628 62475
rect 1618 62389 1628 62445
rect 104 62359 130 62389
rect 1580 62359 1628 62389
rect 1618 62303 1628 62359
rect 104 62273 130 62303
rect 1580 62273 1628 62303
rect 1618 62217 1628 62273
rect 104 62187 130 62217
rect 1580 62187 1628 62217
rect 1618 62131 1628 62187
rect 104 62101 130 62131
rect 1580 62101 1628 62131
rect 1618 62045 1628 62101
rect 104 62015 130 62045
rect 1580 62015 1628 62045
rect 1618 61959 1628 62015
rect 104 61929 130 61959
rect 1580 61929 1628 61959
rect 1618 61873 1628 61929
rect 104 61843 130 61873
rect 1580 61843 1628 61873
rect 1618 61787 1628 61843
rect 104 61757 130 61787
rect 1580 61757 1628 61787
rect 1618 61701 1628 61757
rect 104 61671 130 61701
rect 1580 61671 1628 61701
rect 1618 61615 1628 61671
rect 104 61585 130 61615
rect 1580 61585 1628 61615
rect 1618 61529 1628 61585
rect 104 61499 130 61529
rect 1580 61499 1628 61529
rect 1618 61443 1628 61499
rect 104 61413 130 61443
rect 1580 61413 1628 61443
rect 1618 61357 1628 61413
rect 104 61327 130 61357
rect 1580 61327 1628 61357
rect 1618 61271 1628 61327
rect 104 61241 130 61271
rect 1580 61241 1628 61271
rect 1618 61185 1628 61241
rect 104 61155 130 61185
rect 1580 61155 1628 61185
rect 1618 61099 1628 61155
rect 104 61069 130 61099
rect 1580 61069 1628 61099
rect 1618 61013 1628 61069
rect 104 60983 130 61013
rect 1580 60983 1628 61013
rect 1618 60927 1628 60983
rect 104 60897 130 60927
rect 1580 60897 1628 60927
rect 1618 60841 1628 60897
rect 104 60811 130 60841
rect 1580 60811 1628 60841
rect 1618 60755 1628 60811
rect 104 60725 130 60755
rect 1580 60725 1628 60755
rect 1618 60669 1628 60725
rect 104 60639 130 60669
rect 1580 60639 1628 60669
rect 1618 60583 1628 60639
rect 104 60553 130 60583
rect 1580 60553 1628 60583
rect 1618 60497 1628 60553
rect 104 60467 130 60497
rect 1580 60467 1628 60497
rect 1618 60411 1628 60467
rect 104 60381 130 60411
rect 1580 60381 1628 60411
rect 1618 60325 1628 60381
rect 104 60295 130 60325
rect 1580 60295 1628 60325
rect 1618 60239 1628 60295
rect 104 60209 130 60239
rect 1580 60209 1628 60239
rect 1618 60153 1628 60209
rect 104 60123 130 60153
rect 1580 60123 1628 60153
rect 1618 60067 1628 60123
rect 104 60037 130 60067
rect 1580 60037 1628 60067
rect 1618 59981 1628 60037
rect 104 59951 130 59981
rect 1580 59951 1628 59981
rect 1618 59895 1628 59951
rect 104 59865 130 59895
rect 1580 59865 1628 59895
rect 1618 59809 1628 59865
rect 104 59779 130 59809
rect 1580 59779 1628 59809
rect 1618 59723 1628 59779
rect 104 59693 130 59723
rect 1580 59693 1628 59723
rect 1618 59637 1628 59693
rect 104 59607 130 59637
rect 1580 59607 1628 59637
rect 1618 59551 1628 59607
rect 104 59521 130 59551
rect 1580 59521 1628 59551
rect 1618 59465 1628 59521
rect 104 59435 130 59465
rect 1580 59435 1628 59465
rect 1618 59379 1628 59435
rect 104 59349 130 59379
rect 1580 59349 1628 59379
rect 1618 59293 1628 59349
rect 104 59263 130 59293
rect 1580 59263 1628 59293
rect 1618 59207 1628 59263
rect 104 59177 130 59207
rect 1580 59177 1628 59207
rect 1618 59121 1628 59177
rect 104 59091 130 59121
rect 1580 59091 1628 59121
rect 1618 59035 1628 59091
rect 104 59005 130 59035
rect 1580 59005 1628 59035
rect 1618 58949 1628 59005
rect 104 58919 130 58949
rect 1580 58919 1628 58949
rect 1618 58863 1628 58919
rect 104 58833 130 58863
rect 1580 58833 1628 58863
rect 1618 58777 1628 58833
rect 104 58747 130 58777
rect 1580 58747 1628 58777
rect 1618 58691 1628 58747
rect 104 58661 130 58691
rect 1580 58661 1628 58691
rect 1618 58605 1628 58661
rect 104 58575 130 58605
rect 1580 58575 1628 58605
rect 1618 58519 1628 58575
rect 104 58489 130 58519
rect 1580 58489 1628 58519
rect 1618 58433 1628 58489
rect 104 58403 130 58433
rect 1580 58403 1628 58433
rect 1618 58347 1628 58403
rect 104 58317 130 58347
rect 1580 58317 1628 58347
rect 1618 58261 1628 58317
rect 104 58231 130 58261
rect 1580 58231 1628 58261
rect 1618 58175 1628 58231
rect 104 58145 130 58175
rect 1580 58145 1628 58175
rect 1618 58089 1628 58145
rect 104 58059 130 58089
rect 1580 58059 1628 58089
rect 1618 58003 1628 58059
rect 104 57973 130 58003
rect 1580 57973 1628 58003
rect 1618 57917 1628 57973
rect 104 57887 130 57917
rect 1580 57887 1628 57917
rect 1618 57831 1628 57887
rect 104 57801 130 57831
rect 1580 57801 1628 57831
rect 1618 57745 1628 57801
rect 104 57715 130 57745
rect 1580 57715 1628 57745
rect 1618 57659 1628 57715
rect 104 57629 130 57659
rect 1580 57629 1628 57659
rect 1618 57573 1628 57629
rect 104 57543 130 57573
rect 1580 57543 1628 57573
rect 1618 57487 1628 57543
rect 104 57457 130 57487
rect 1580 57457 1628 57487
rect 1618 57401 1628 57457
rect 104 57371 130 57401
rect 1580 57371 1628 57401
rect 1618 57315 1628 57371
rect 104 57285 130 57315
rect 1580 57285 1628 57315
rect 1618 57229 1628 57285
rect 104 57199 130 57229
rect 1580 57199 1628 57229
rect 1618 57143 1628 57199
rect 104 57113 130 57143
rect 1580 57113 1628 57143
rect 1618 57057 1628 57113
rect 104 57027 130 57057
rect 1580 57027 1628 57057
rect 1618 56971 1628 57027
rect 104 56941 130 56971
rect 1580 56941 1628 56971
rect 1618 56885 1628 56941
rect 104 56855 130 56885
rect 1580 56855 1628 56885
rect 1618 56799 1628 56855
rect 104 56769 130 56799
rect 1580 56769 1628 56799
rect 1618 56713 1628 56769
rect 104 56683 130 56713
rect 1580 56683 1628 56713
rect 1618 56627 1628 56683
rect 104 56597 130 56627
rect 1580 56597 1628 56627
rect 1618 56541 1628 56597
rect 104 56511 130 56541
rect 1580 56511 1628 56541
rect 1618 56455 1628 56511
rect 104 56425 130 56455
rect 1580 56425 1628 56455
rect 1618 56369 1628 56425
rect 104 56339 130 56369
rect 1580 56339 1628 56369
rect 1618 56283 1628 56339
rect 104 56253 130 56283
rect 1580 56253 1628 56283
rect 1618 56197 1628 56253
rect 104 56167 130 56197
rect 1580 56167 1628 56197
rect 1618 56111 1628 56167
rect 104 56081 130 56111
rect 1580 56081 1628 56111
rect 1618 56025 1628 56081
rect 104 55995 130 56025
rect 1580 55995 1628 56025
rect 1618 55939 1628 55995
rect 104 55909 130 55939
rect 1580 55909 1628 55939
rect 1618 55853 1628 55909
rect 104 55823 130 55853
rect 1580 55823 1628 55853
rect 1618 55767 1628 55823
rect 104 55737 130 55767
rect 1580 55737 1628 55767
rect 1618 55681 1628 55737
rect 104 55651 130 55681
rect 1580 55651 1628 55681
rect 1618 55595 1628 55651
rect 104 55565 130 55595
rect 1580 55565 1628 55595
rect 1618 55509 1628 55565
rect 104 55479 130 55509
rect 1580 55479 1628 55509
rect 1618 55423 1628 55479
rect 104 55393 130 55423
rect 1580 55393 1628 55423
rect 1618 55337 1628 55393
rect 104 55307 130 55337
rect 1580 55307 1628 55337
rect 1618 55251 1628 55307
rect 104 55221 130 55251
rect 1580 55221 1628 55251
rect 1618 55165 1628 55221
rect 104 55135 130 55165
rect 1580 55135 1628 55165
rect 1618 55079 1628 55135
rect 104 55049 130 55079
rect 1580 55049 1628 55079
rect 1618 54993 1628 55049
rect 104 54963 130 54993
rect 1580 54963 1628 54993
rect 1618 54907 1628 54963
rect 104 54877 130 54907
rect 1580 54877 1628 54907
rect 1618 54821 1628 54877
rect 104 54791 130 54821
rect 1580 54791 1628 54821
rect 1618 54735 1628 54791
rect 104 54705 130 54735
rect 1580 54705 1628 54735
rect 1618 54649 1628 54705
rect 104 54619 130 54649
rect 1580 54619 1628 54649
rect 1618 54563 1628 54619
rect 104 54533 130 54563
rect 1580 54533 1628 54563
rect 1618 54477 1628 54533
rect 104 54447 130 54477
rect 1580 54447 1628 54477
rect 1618 54391 1628 54447
rect 104 54361 130 54391
rect 1580 54361 1628 54391
rect 1618 54305 1628 54361
rect 104 54275 130 54305
rect 1580 54275 1628 54305
rect 1618 54219 1628 54275
rect 104 54189 130 54219
rect 1580 54189 1628 54219
rect 1618 54133 1628 54189
rect 104 54103 130 54133
rect 1580 54103 1628 54133
rect 1618 54047 1628 54103
rect 104 54017 130 54047
rect 1580 54017 1628 54047
rect 1618 53961 1628 54017
rect 104 53931 130 53961
rect 1580 53931 1628 53961
rect 1618 53875 1628 53931
rect 104 53845 130 53875
rect 1580 53845 1628 53875
rect 1618 53789 1628 53845
rect 104 53759 130 53789
rect 1580 53759 1628 53789
rect 1618 53703 1628 53759
rect 104 53673 130 53703
rect 1580 53673 1628 53703
rect 1618 53617 1628 53673
rect 104 53587 130 53617
rect 1580 53587 1628 53617
rect 1618 53531 1628 53587
rect 104 53501 130 53531
rect 1580 53501 1628 53531
rect 1618 53445 1628 53501
rect 104 53415 130 53445
rect 1580 53415 1628 53445
rect 1618 53359 1628 53415
rect 104 53329 130 53359
rect 1580 53329 1628 53359
rect 1618 53273 1628 53329
rect 104 53243 130 53273
rect 1580 53243 1628 53273
rect 1618 53187 1628 53243
rect 104 53157 130 53187
rect 1580 53157 1628 53187
rect 1618 53101 1628 53157
rect 104 53071 130 53101
rect 1580 53071 1628 53101
rect 1618 53015 1628 53071
rect 104 52985 130 53015
rect 1580 52985 1628 53015
rect 1618 52929 1628 52985
rect 104 52899 130 52929
rect 1580 52899 1628 52929
rect 1618 52843 1628 52899
rect 104 52813 130 52843
rect 1580 52813 1628 52843
rect 1618 52757 1628 52813
rect 104 52727 130 52757
rect 1580 52727 1628 52757
rect 1618 52671 1628 52727
rect 104 52641 130 52671
rect 1580 52641 1628 52671
rect 1618 52585 1628 52641
rect 104 52555 130 52585
rect 1580 52555 1628 52585
rect 1618 52499 1628 52555
rect 104 52469 130 52499
rect 1580 52469 1628 52499
rect 1618 52413 1628 52469
rect 104 52383 130 52413
rect 1580 52383 1628 52413
rect 1618 52327 1628 52383
rect 104 52297 130 52327
rect 1580 52297 1628 52327
rect 1618 52241 1628 52297
rect 104 52211 130 52241
rect 1580 52211 1628 52241
rect 1618 52155 1628 52211
rect 104 52125 130 52155
rect 1580 52125 1628 52155
rect 1618 52069 1628 52125
rect 104 52039 130 52069
rect 1580 52039 1628 52069
rect 1618 51983 1628 52039
rect 104 51953 130 51983
rect 1580 51953 1628 51983
rect 1618 51897 1628 51953
rect 104 51867 130 51897
rect 1580 51867 1628 51897
rect 1618 51811 1628 51867
rect 104 51781 130 51811
rect 1580 51781 1628 51811
rect 1618 51725 1628 51781
rect 104 51695 130 51725
rect 1580 51695 1628 51725
rect 1618 51639 1628 51695
rect 104 51609 130 51639
rect 1580 51609 1628 51639
rect 1618 51553 1628 51609
rect 104 51523 130 51553
rect 1580 51523 1628 51553
rect 1618 51467 1628 51523
rect 104 51437 130 51467
rect 1580 51437 1628 51467
rect 1618 51381 1628 51437
rect 104 51351 130 51381
rect 1580 51351 1628 51381
rect 1618 51295 1628 51351
rect 104 51265 130 51295
rect 1580 51265 1628 51295
rect 1618 51209 1628 51265
rect 104 51179 130 51209
rect 1580 51179 1628 51209
rect 1618 51123 1628 51179
rect 104 51093 130 51123
rect 1580 51093 1628 51123
rect 1618 51037 1628 51093
rect 104 51007 130 51037
rect 1580 51007 1628 51037
rect 1618 50951 1628 51007
rect 104 50921 130 50951
rect 1580 50921 1628 50951
rect 1618 50865 1628 50921
rect 104 50835 130 50865
rect 1580 50835 1628 50865
rect 1618 50779 1628 50835
rect 104 50749 130 50779
rect 1580 50749 1628 50779
rect 1618 50693 1628 50749
rect 104 50663 130 50693
rect 1580 50663 1628 50693
rect 1618 50607 1628 50663
rect 104 50577 130 50607
rect 1580 50577 1628 50607
rect 1618 50521 1628 50577
rect 104 50491 130 50521
rect 1580 50491 1628 50521
rect 1618 50435 1628 50491
rect 104 50405 130 50435
rect 1580 50405 1628 50435
rect 1618 50349 1628 50405
rect 104 50319 130 50349
rect 1580 50319 1628 50349
rect 1618 50263 1628 50319
rect 104 50233 130 50263
rect 1580 50233 1628 50263
rect 1618 50177 1628 50233
rect 104 50147 130 50177
rect 1580 50147 1628 50177
rect 1618 50091 1628 50147
rect 104 50061 130 50091
rect 1580 50061 1628 50091
rect 1618 50005 1628 50061
rect 104 49975 130 50005
rect 1580 49975 1628 50005
rect 1618 49919 1628 49975
rect 104 49889 130 49919
rect 1580 49889 1628 49919
rect 1618 49833 1628 49889
rect 104 49803 130 49833
rect 1580 49803 1628 49833
rect 1618 49747 1628 49803
rect 104 49717 130 49747
rect 1580 49717 1628 49747
rect 1618 49661 1628 49717
rect 104 49631 130 49661
rect 1580 49631 1628 49661
rect 1618 49575 1628 49631
rect 104 49545 130 49575
rect 1580 49545 1628 49575
rect 1618 49489 1628 49545
rect 104 49459 130 49489
rect 1580 49459 1628 49489
rect 1618 49403 1628 49459
rect 104 49373 130 49403
rect 1580 49373 1628 49403
rect 1618 49317 1628 49373
rect 104 49287 130 49317
rect 1580 49287 1628 49317
rect 1618 49231 1628 49287
rect 104 49201 130 49231
rect 1580 49201 1628 49231
rect 1618 49145 1628 49201
rect 104 49115 130 49145
rect 1580 49115 1628 49145
rect 1618 49059 1628 49115
rect 104 49029 130 49059
rect 1580 49029 1628 49059
rect 1618 48973 1628 49029
rect 104 48943 130 48973
rect 1580 48943 1628 48973
rect 1618 48887 1628 48943
rect 104 48857 130 48887
rect 1580 48857 1628 48887
rect 1618 48801 1628 48857
rect 104 48771 130 48801
rect 1580 48771 1628 48801
rect 1618 48715 1628 48771
rect 104 48685 130 48715
rect 1580 48685 1628 48715
rect 1618 48629 1628 48685
rect 104 48599 130 48629
rect 1580 48599 1628 48629
rect 1618 48543 1628 48599
rect 104 48513 130 48543
rect 1580 48513 1628 48543
rect 1618 48457 1628 48513
rect 104 48427 130 48457
rect 1580 48427 1628 48457
rect 1618 48371 1628 48427
rect 104 48341 130 48371
rect 1580 48341 1628 48371
rect 1618 48285 1628 48341
rect 104 48255 130 48285
rect 1580 48255 1628 48285
rect 1618 48199 1628 48255
rect 104 48169 130 48199
rect 1580 48169 1628 48199
rect 1618 48113 1628 48169
rect 104 48083 130 48113
rect 1580 48083 1628 48113
rect 1618 48027 1628 48083
rect 104 47997 130 48027
rect 1580 47997 1628 48027
rect 1618 47941 1628 47997
rect 104 47911 130 47941
rect 1580 47911 1628 47941
rect 1618 47855 1628 47911
rect 104 47825 130 47855
rect 1580 47825 1628 47855
rect 1618 47769 1628 47825
rect 104 47739 130 47769
rect 1580 47739 1628 47769
rect 1618 47683 1628 47739
rect 104 47653 130 47683
rect 1580 47653 1628 47683
rect 1618 47597 1628 47653
rect 104 47567 130 47597
rect 1580 47567 1628 47597
rect 1618 47511 1628 47567
rect 104 47481 130 47511
rect 1580 47481 1628 47511
rect 1618 47425 1628 47481
rect 104 47395 130 47425
rect 1580 47395 1628 47425
rect 1618 47339 1628 47395
rect 104 47309 130 47339
rect 1580 47309 1628 47339
rect 1618 47253 1628 47309
rect 104 47223 130 47253
rect 1580 47223 1628 47253
rect 1618 47167 1628 47223
rect 104 47137 130 47167
rect 1580 47137 1628 47167
rect 1618 47081 1628 47137
rect 104 47051 130 47081
rect 1580 47051 1628 47081
rect 1618 46995 1628 47051
rect 104 46965 130 46995
rect 1580 46965 1628 46995
rect 1618 46909 1628 46965
rect 104 46879 130 46909
rect 1580 46879 1628 46909
rect 1618 46823 1628 46879
rect 104 46793 130 46823
rect 1580 46793 1628 46823
rect 1618 46737 1628 46793
rect 104 46707 130 46737
rect 1580 46707 1628 46737
rect 1618 46651 1628 46707
rect 104 46621 130 46651
rect 1580 46621 1628 46651
rect 1618 46565 1628 46621
rect 104 46535 130 46565
rect 1580 46535 1628 46565
rect 1618 46479 1628 46535
rect 104 46449 130 46479
rect 1580 46449 1628 46479
rect 1618 46393 1628 46449
rect 104 46363 130 46393
rect 1580 46363 1628 46393
rect 1618 46307 1628 46363
rect 104 46277 130 46307
rect 1580 46277 1628 46307
rect 1618 46221 1628 46277
rect 104 46191 130 46221
rect 1580 46191 1628 46221
rect 1618 46135 1628 46191
rect 104 46105 130 46135
rect 1580 46105 1628 46135
rect 1618 46049 1628 46105
rect 104 46019 130 46049
rect 1580 46019 1628 46049
rect 1618 45963 1628 46019
rect 104 45933 130 45963
rect 1580 45933 1628 45963
rect 1618 45877 1628 45933
rect 104 45847 130 45877
rect 1580 45847 1628 45877
rect 1618 45791 1628 45847
rect 104 45761 130 45791
rect 1580 45761 1628 45791
rect 1618 45705 1628 45761
rect 104 45675 130 45705
rect 1580 45675 1628 45705
rect 1618 45619 1628 45675
rect 104 45589 130 45619
rect 1580 45589 1628 45619
rect 1618 45533 1628 45589
rect 104 45503 130 45533
rect 1580 45503 1628 45533
rect 1618 45447 1628 45503
rect 104 45417 130 45447
rect 1580 45417 1628 45447
rect 1618 45361 1628 45417
rect 104 45331 130 45361
rect 1580 45331 1628 45361
rect 1618 45275 1628 45331
rect 104 45245 130 45275
rect 1580 45245 1628 45275
rect 1618 45189 1628 45245
rect 104 45159 130 45189
rect 1580 45159 1628 45189
rect 1618 45103 1628 45159
rect 104 45073 130 45103
rect 1580 45073 1628 45103
rect 1618 45017 1628 45073
rect 104 44987 130 45017
rect 1580 44987 1628 45017
rect 1618 44931 1628 44987
rect 104 44901 130 44931
rect 1580 44901 1628 44931
rect 1618 44845 1628 44901
rect 104 44815 130 44845
rect 1580 44815 1628 44845
rect 1618 44759 1628 44815
rect 104 44729 130 44759
rect 1580 44729 1628 44759
rect 1618 44673 1628 44729
rect 104 44643 130 44673
rect 1580 44643 1628 44673
rect 1618 44587 1628 44643
rect 104 44557 130 44587
rect 1580 44557 1628 44587
rect 1618 44501 1628 44557
rect 104 44471 130 44501
rect 1580 44471 1628 44501
rect 1618 44415 1628 44471
rect 104 44385 130 44415
rect 1580 44385 1628 44415
rect 1618 44329 1628 44385
rect 104 44299 130 44329
rect 1580 44299 1628 44329
rect 1618 44243 1628 44299
rect 104 44213 130 44243
rect 1580 44213 1628 44243
rect 1618 44157 1628 44213
rect 104 44127 130 44157
rect 1580 44127 1628 44157
rect 1618 44071 1628 44127
rect 104 44041 130 44071
rect 1580 44041 1628 44071
rect 1618 43985 1628 44041
rect 104 43955 130 43985
rect 1580 43955 1628 43985
rect 1618 43899 1628 43955
rect 104 43869 130 43899
rect 1580 43869 1628 43899
rect 1618 43813 1628 43869
rect 104 43783 130 43813
rect 1580 43783 1628 43813
rect 1618 43727 1628 43783
rect 104 43697 130 43727
rect 1580 43697 1628 43727
rect 1618 43641 1628 43697
rect 104 43611 130 43641
rect 1580 43611 1628 43641
rect 1618 43555 1628 43611
rect 104 43525 130 43555
rect 1580 43525 1628 43555
rect 1618 43469 1628 43525
rect 104 43439 130 43469
rect 1580 43439 1628 43469
rect 1618 43383 1628 43439
rect 104 43353 130 43383
rect 1580 43353 1628 43383
rect 1618 43297 1628 43353
rect 104 43267 130 43297
rect 1580 43267 1628 43297
rect 1618 43211 1628 43267
rect 104 43181 130 43211
rect 1580 43181 1628 43211
rect 1618 43125 1628 43181
rect 104 43095 130 43125
rect 1580 43095 1628 43125
rect 1618 43039 1628 43095
rect 104 43009 130 43039
rect 1580 43009 1628 43039
rect 1618 42953 1628 43009
rect 104 42923 130 42953
rect 1580 42923 1628 42953
rect 1618 42867 1628 42923
rect 104 42837 130 42867
rect 1580 42837 1628 42867
rect 1618 42781 1628 42837
rect 104 42751 130 42781
rect 1580 42751 1628 42781
rect 1618 42695 1628 42751
rect 104 42665 130 42695
rect 1580 42665 1628 42695
rect 1618 42609 1628 42665
rect 104 42579 130 42609
rect 1580 42579 1628 42609
rect 1618 42523 1628 42579
rect 104 42493 130 42523
rect 1580 42493 1628 42523
rect 1618 42437 1628 42493
rect 104 42407 130 42437
rect 1580 42407 1628 42437
rect 1618 42351 1628 42407
rect 104 42321 130 42351
rect 1580 42321 1628 42351
rect 1618 42265 1628 42321
rect 104 42235 130 42265
rect 1580 42235 1628 42265
rect 1618 42179 1628 42235
rect 104 42149 130 42179
rect 1580 42149 1628 42179
rect 1618 42093 1628 42149
rect 104 42063 130 42093
rect 1580 42063 1628 42093
rect 1618 42007 1628 42063
rect 104 41977 130 42007
rect 1580 41977 1628 42007
rect 1618 41921 1628 41977
rect 104 41891 130 41921
rect 1580 41891 1628 41921
rect 1618 41835 1628 41891
rect 104 41805 130 41835
rect 1580 41805 1628 41835
rect 1618 41749 1628 41805
rect 104 41719 130 41749
rect 1580 41719 1628 41749
rect 1618 41663 1628 41719
rect 104 41633 130 41663
rect 1580 41633 1628 41663
rect 1618 41577 1628 41633
rect 104 41547 130 41577
rect 1580 41547 1628 41577
rect 1618 41491 1628 41547
rect 104 41461 130 41491
rect 1580 41461 1628 41491
rect 1618 41405 1628 41461
rect 104 41375 130 41405
rect 1580 41375 1628 41405
rect 1618 41319 1628 41375
rect 104 41289 130 41319
rect 1580 41289 1628 41319
rect 1618 41233 1628 41289
rect 104 41203 130 41233
rect 1580 41203 1628 41233
rect 1618 41147 1628 41203
rect 104 41117 130 41147
rect 1580 41117 1628 41147
rect 1618 41061 1628 41117
rect 104 41031 130 41061
rect 1580 41031 1628 41061
rect 1618 40975 1628 41031
rect 104 40945 130 40975
rect 1580 40945 1628 40975
rect 1618 40889 1628 40945
rect 104 40859 130 40889
rect 1580 40859 1628 40889
rect 1618 40803 1628 40859
rect 104 40773 130 40803
rect 1580 40773 1628 40803
rect 1618 40717 1628 40773
rect 104 40687 130 40717
rect 1580 40687 1628 40717
rect 1618 40631 1628 40687
rect 104 40601 130 40631
rect 1580 40601 1628 40631
rect 1618 40545 1628 40601
rect 104 40515 130 40545
rect 1580 40515 1628 40545
rect 1618 40459 1628 40515
rect 104 40429 130 40459
rect 1580 40429 1628 40459
rect 1618 40373 1628 40429
rect 104 40343 130 40373
rect 1580 40343 1628 40373
rect 1618 40287 1628 40343
rect 104 40257 130 40287
rect 1580 40257 1628 40287
rect 1618 40201 1628 40257
rect 104 40171 130 40201
rect 1580 40171 1628 40201
rect 1618 40115 1628 40171
rect 104 40085 130 40115
rect 1580 40085 1628 40115
rect 1618 40029 1628 40085
rect 104 39999 130 40029
rect 1580 39999 1628 40029
rect 1618 39943 1628 39999
rect 104 39913 130 39943
rect 1580 39913 1628 39943
rect 1618 39857 1628 39913
rect 104 39827 130 39857
rect 1580 39827 1628 39857
rect 1618 39771 1628 39827
rect 104 39741 130 39771
rect 1580 39741 1628 39771
rect 1618 39685 1628 39741
rect 104 39655 130 39685
rect 1580 39655 1628 39685
rect 1618 39599 1628 39655
rect 104 39569 130 39599
rect 1580 39569 1628 39599
rect 1618 39513 1628 39569
rect 104 39483 130 39513
rect 1580 39483 1628 39513
rect 1618 39427 1628 39483
rect 104 39397 130 39427
rect 1580 39397 1628 39427
rect 1618 39341 1628 39397
rect 104 39311 130 39341
rect 1580 39311 1628 39341
rect 1618 39255 1628 39311
rect 104 39225 130 39255
rect 1580 39225 1628 39255
rect 1618 39169 1628 39225
rect 104 39139 130 39169
rect 1580 39139 1628 39169
rect 1618 39083 1628 39139
rect 104 39053 130 39083
rect 1580 39053 1628 39083
rect 1618 38997 1628 39053
rect 104 38967 130 38997
rect 1580 38967 1628 38997
rect 1618 38911 1628 38967
rect 104 38881 130 38911
rect 1580 38881 1628 38911
rect 1618 38825 1628 38881
rect 104 38795 130 38825
rect 1580 38795 1628 38825
rect 1618 38739 1628 38795
rect 104 38709 130 38739
rect 1580 38709 1628 38739
rect 1618 38653 1628 38709
rect 104 38623 130 38653
rect 1580 38623 1628 38653
rect 1618 38567 1628 38623
rect 104 38537 130 38567
rect 1580 38537 1628 38567
rect 1618 38481 1628 38537
rect 104 38451 130 38481
rect 1580 38451 1628 38481
rect 1618 38395 1628 38451
rect 104 38365 130 38395
rect 1580 38365 1628 38395
rect 1618 38309 1628 38365
rect 104 38279 130 38309
rect 1580 38279 1628 38309
rect 1618 38223 1628 38279
rect 104 38193 130 38223
rect 1580 38193 1628 38223
rect 1618 38137 1628 38193
rect 104 38107 130 38137
rect 1580 38107 1628 38137
rect 1618 38051 1628 38107
rect 104 38021 130 38051
rect 1580 38021 1628 38051
rect 1618 37965 1628 38021
rect 104 37935 130 37965
rect 1580 37935 1628 37965
rect 1618 37879 1628 37935
rect 104 37849 130 37879
rect 1580 37849 1628 37879
rect 1618 37793 1628 37849
rect 104 37763 130 37793
rect 1580 37763 1628 37793
rect 1618 37707 1628 37763
rect 104 37677 130 37707
rect 1580 37677 1628 37707
rect 1618 37621 1628 37677
rect 104 37591 130 37621
rect 1580 37591 1628 37621
rect 1618 37535 1628 37591
rect 104 37505 130 37535
rect 1580 37505 1628 37535
rect 1618 37449 1628 37505
rect 104 37419 130 37449
rect 1580 37419 1628 37449
rect 1618 37363 1628 37419
rect 104 37333 130 37363
rect 1580 37333 1628 37363
rect 1618 37277 1628 37333
rect 104 37247 130 37277
rect 1580 37247 1628 37277
rect 1618 37191 1628 37247
rect 104 37161 130 37191
rect 1580 37161 1628 37191
rect 1618 37105 1628 37161
rect 104 37075 130 37105
rect 1580 37075 1628 37105
rect 1618 37019 1628 37075
rect 104 36989 130 37019
rect 1580 36989 1628 37019
rect 1618 36933 1628 36989
rect 104 36903 130 36933
rect 1580 36903 1628 36933
rect 1618 36847 1628 36903
rect 104 36817 130 36847
rect 1580 36817 1628 36847
rect 1618 36761 1628 36817
rect 104 36731 130 36761
rect 1580 36731 1628 36761
rect 1618 36675 1628 36731
rect 104 36645 130 36675
rect 1580 36645 1628 36675
rect 1618 36589 1628 36645
rect 104 36559 130 36589
rect 1580 36559 1628 36589
rect 1618 36503 1628 36559
rect 104 36473 130 36503
rect 1580 36473 1628 36503
rect 1618 36417 1628 36473
rect 104 36387 130 36417
rect 1580 36387 1628 36417
rect 1618 36331 1628 36387
rect 104 36301 130 36331
rect 1580 36301 1628 36331
rect 1618 36245 1628 36301
rect 104 36215 130 36245
rect 1580 36215 1628 36245
rect 1618 36159 1628 36215
rect 104 36129 130 36159
rect 1580 36129 1628 36159
rect 1618 36073 1628 36129
rect 104 36043 130 36073
rect 1580 36043 1628 36073
rect 1618 35987 1628 36043
rect 104 35957 130 35987
rect 1580 35957 1628 35987
rect 1618 35901 1628 35957
rect 104 35871 130 35901
rect 1580 35871 1628 35901
rect 1618 35815 1628 35871
rect 104 35785 130 35815
rect 1580 35785 1628 35815
rect 1618 35729 1628 35785
rect 104 35699 130 35729
rect 1580 35699 1628 35729
rect 1618 35643 1628 35699
rect 104 35613 130 35643
rect 1580 35613 1628 35643
rect 1618 35557 1628 35613
rect 104 35527 130 35557
rect 1580 35527 1628 35557
rect 1618 35471 1628 35527
rect 104 35441 130 35471
rect 1580 35441 1628 35471
rect 1618 35385 1628 35441
rect 104 35355 130 35385
rect 1580 35355 1628 35385
rect 1618 35299 1628 35355
rect 104 35269 130 35299
rect 1580 35269 1628 35299
rect 1618 35213 1628 35269
rect 104 35183 130 35213
rect 1580 35183 1628 35213
rect 1618 35127 1628 35183
rect 104 35097 130 35127
rect 1580 35097 1628 35127
rect 1618 35041 1628 35097
rect 104 35011 130 35041
rect 1580 35011 1628 35041
rect 1618 34955 1628 35011
rect 104 34925 130 34955
rect 1580 34925 1628 34955
rect 1618 34869 1628 34925
rect 104 34839 130 34869
rect 1580 34839 1628 34869
rect 1618 34783 1628 34839
rect 104 34753 130 34783
rect 1580 34753 1628 34783
rect 1618 34697 1628 34753
rect 104 34667 130 34697
rect 1580 34667 1628 34697
rect 1618 34611 1628 34667
rect 104 34581 130 34611
rect 1580 34581 1628 34611
rect 1618 34525 1628 34581
rect 104 34495 130 34525
rect 1580 34495 1628 34525
rect 1618 34439 1628 34495
rect 104 34409 130 34439
rect 1580 34409 1628 34439
rect 1618 34353 1628 34409
rect 104 34323 130 34353
rect 1580 34323 1628 34353
rect 1618 34267 1628 34323
rect 104 34237 130 34267
rect 1580 34237 1628 34267
rect 1618 34181 1628 34237
rect 104 34151 130 34181
rect 1580 34151 1628 34181
rect 1618 34095 1628 34151
rect 104 34065 130 34095
rect 1580 34065 1628 34095
rect 1618 34009 1628 34065
rect 104 33979 130 34009
rect 1580 33979 1628 34009
rect 1618 33923 1628 33979
rect 104 33893 130 33923
rect 1580 33893 1628 33923
rect 1618 33837 1628 33893
rect 104 33807 130 33837
rect 1580 33807 1628 33837
rect 1618 33751 1628 33807
rect 104 33721 130 33751
rect 1580 33721 1628 33751
rect 1618 33665 1628 33721
rect 104 33635 130 33665
rect 1580 33635 1628 33665
rect 1618 33579 1628 33635
rect 104 33549 130 33579
rect 1580 33549 1628 33579
rect 1618 33493 1628 33549
rect 104 33463 130 33493
rect 1580 33463 1628 33493
rect 1618 33407 1628 33463
rect 104 33377 130 33407
rect 1580 33377 1628 33407
rect 1618 33321 1628 33377
rect 104 33291 130 33321
rect 1580 33291 1628 33321
rect 1618 33235 1628 33291
rect 104 33205 130 33235
rect 1580 33205 1628 33235
rect 1618 33149 1628 33205
rect 104 33119 130 33149
rect 1580 33119 1628 33149
rect 1618 33063 1628 33119
rect 104 33033 130 33063
rect 1580 33033 1628 33063
rect 1618 32977 1628 33033
rect 104 32947 130 32977
rect 1580 32947 1628 32977
rect 1618 32891 1628 32947
rect 104 32861 130 32891
rect 1580 32861 1628 32891
rect 1618 32805 1628 32861
rect 104 32775 130 32805
rect 1580 32775 1628 32805
rect 1618 32719 1628 32775
rect 104 32689 130 32719
rect 1580 32689 1628 32719
rect 1618 32633 1628 32689
rect 104 32603 130 32633
rect 1580 32603 1628 32633
rect 1618 32547 1628 32603
rect 104 32517 130 32547
rect 1580 32517 1628 32547
rect 1618 32461 1628 32517
rect 104 32431 130 32461
rect 1580 32431 1628 32461
rect 1618 32375 1628 32431
rect 104 32345 130 32375
rect 1580 32345 1628 32375
rect 1618 32289 1628 32345
rect 104 32259 130 32289
rect 1580 32259 1628 32289
rect 1618 32203 1628 32259
rect 104 32173 130 32203
rect 1580 32173 1628 32203
rect 1618 32117 1628 32173
rect 104 32087 130 32117
rect 1580 32087 1628 32117
rect 1618 32031 1628 32087
rect 104 32001 130 32031
rect 1580 32001 1628 32031
rect 1618 31945 1628 32001
rect 104 31915 130 31945
rect 1580 31915 1628 31945
rect 1618 31859 1628 31915
rect 104 31829 130 31859
rect 1580 31829 1628 31859
rect 1618 31773 1628 31829
rect 104 31743 130 31773
rect 1580 31743 1628 31773
rect 1618 31687 1628 31743
rect 104 31657 130 31687
rect 1580 31657 1628 31687
rect 1618 31601 1628 31657
rect 104 31571 130 31601
rect 1580 31571 1628 31601
rect 1618 31515 1628 31571
rect 104 31485 130 31515
rect 1580 31485 1628 31515
rect 1618 31429 1628 31485
rect 104 31399 130 31429
rect 1580 31399 1628 31429
rect 1618 31343 1628 31399
rect 104 31313 130 31343
rect 1580 31313 1628 31343
rect 1618 31257 1628 31313
rect 104 31227 130 31257
rect 1580 31227 1628 31257
rect 1618 31171 1628 31227
rect 104 31141 130 31171
rect 1580 31141 1628 31171
rect 1618 31085 1628 31141
rect 104 31055 130 31085
rect 1580 31055 1628 31085
rect 1618 30999 1628 31055
rect 104 30969 130 30999
rect 1580 30969 1628 30999
rect 1618 30913 1628 30969
rect 104 30883 130 30913
rect 1580 30883 1628 30913
rect 1618 30827 1628 30883
rect 104 30797 130 30827
rect 1580 30797 1628 30827
rect 1618 30741 1628 30797
rect 104 30711 130 30741
rect 1580 30711 1628 30741
rect 1618 30655 1628 30711
rect 104 30625 130 30655
rect 1580 30625 1628 30655
rect 1618 30569 1628 30625
rect 104 30539 130 30569
rect 1580 30539 1628 30569
rect 1618 30483 1628 30539
rect 104 30453 130 30483
rect 1580 30453 1628 30483
rect 1618 30397 1628 30453
rect 104 30367 130 30397
rect 1580 30367 1628 30397
rect 1618 30311 1628 30367
rect 104 30281 130 30311
rect 1580 30281 1628 30311
rect 1618 30225 1628 30281
rect 104 30195 130 30225
rect 1580 30195 1628 30225
rect 1618 30139 1628 30195
rect 104 30109 130 30139
rect 1580 30109 1628 30139
rect 1618 30053 1628 30109
rect 104 30023 130 30053
rect 1580 30023 1628 30053
rect 1618 29967 1628 30023
rect 104 29937 130 29967
rect 1580 29937 1628 29967
rect 1618 29881 1628 29937
rect 104 29851 130 29881
rect 1580 29851 1628 29881
rect 1618 29795 1628 29851
rect 104 29765 130 29795
rect 1580 29765 1628 29795
rect 1618 29709 1628 29765
rect 104 29679 130 29709
rect 1580 29679 1628 29709
rect 1618 29623 1628 29679
rect 104 29593 130 29623
rect 1580 29593 1628 29623
rect 1618 29537 1628 29593
rect 104 29507 130 29537
rect 1580 29507 1628 29537
rect 1618 29451 1628 29507
rect 104 29421 130 29451
rect 1580 29421 1628 29451
rect 1618 29365 1628 29421
rect 104 29335 130 29365
rect 1580 29335 1628 29365
rect 1618 29279 1628 29335
rect 104 29249 130 29279
rect 1580 29249 1628 29279
rect 1618 29193 1628 29249
rect 104 29163 130 29193
rect 1580 29163 1628 29193
rect 1618 29107 1628 29163
rect 104 29077 130 29107
rect 1580 29077 1628 29107
rect 1618 29021 1628 29077
rect 104 28991 130 29021
rect 1580 28991 1628 29021
rect 1618 28935 1628 28991
rect 104 28905 130 28935
rect 1580 28905 1628 28935
rect 1618 28849 1628 28905
rect 104 28819 130 28849
rect 1580 28819 1628 28849
rect 1618 28763 1628 28819
rect 104 28733 130 28763
rect 1580 28733 1628 28763
rect 1618 28677 1628 28733
rect 104 28647 130 28677
rect 1580 28647 1628 28677
rect 1618 28591 1628 28647
rect 104 28561 130 28591
rect 1580 28561 1628 28591
rect 1618 28505 1628 28561
rect 104 28475 130 28505
rect 1580 28475 1628 28505
rect 1618 28419 1628 28475
rect 104 28389 130 28419
rect 1580 28389 1628 28419
rect 1618 28333 1628 28389
rect 104 28303 130 28333
rect 1580 28303 1628 28333
rect 1618 28247 1628 28303
rect 104 28217 130 28247
rect 1580 28217 1628 28247
rect 1618 28161 1628 28217
rect 104 28131 130 28161
rect 1580 28131 1628 28161
rect 1618 28075 1628 28131
rect 104 28045 130 28075
rect 1580 28045 1628 28075
rect 1618 27989 1628 28045
rect 104 27959 130 27989
rect 1580 27959 1628 27989
rect 1618 27903 1628 27959
rect 104 27873 130 27903
rect 1580 27873 1628 27903
rect 1618 27817 1628 27873
rect 104 27787 130 27817
rect 1580 27787 1628 27817
rect 1618 27731 1628 27787
rect 104 27701 130 27731
rect 1580 27701 1628 27731
rect 1618 27645 1628 27701
rect 104 27615 130 27645
rect 1580 27615 1628 27645
rect 1618 27559 1628 27615
rect 104 27529 130 27559
rect 1580 27529 1628 27559
rect 1618 27473 1628 27529
rect 104 27443 130 27473
rect 1580 27443 1628 27473
rect 1618 27387 1628 27443
rect 104 27357 130 27387
rect 1580 27357 1628 27387
rect 1618 27301 1628 27357
rect 104 27271 130 27301
rect 1580 27271 1628 27301
rect 1618 27215 1628 27271
rect 104 27185 130 27215
rect 1580 27185 1628 27215
rect 1618 27129 1628 27185
rect 104 27099 130 27129
rect 1580 27099 1628 27129
rect 1618 27043 1628 27099
rect 104 27013 130 27043
rect 1580 27013 1628 27043
rect 1618 26957 1628 27013
rect 104 26927 130 26957
rect 1580 26927 1628 26957
rect 1618 26871 1628 26927
rect 104 26841 130 26871
rect 1580 26841 1628 26871
rect 1618 26785 1628 26841
rect 104 26755 130 26785
rect 1580 26755 1628 26785
rect 1618 26699 1628 26755
rect 104 26669 130 26699
rect 1580 26669 1628 26699
rect 1618 26613 1628 26669
rect 104 26583 130 26613
rect 1580 26583 1628 26613
rect 1618 26527 1628 26583
rect 104 26497 130 26527
rect 1580 26497 1628 26527
rect 1618 26441 1628 26497
rect 104 26411 130 26441
rect 1580 26411 1628 26441
rect 1618 26355 1628 26411
rect 104 26325 130 26355
rect 1580 26325 1628 26355
rect 1618 26269 1628 26325
rect 104 26239 130 26269
rect 1580 26239 1628 26269
rect 1618 26183 1628 26239
rect 104 26153 130 26183
rect 1580 26153 1628 26183
rect 1618 26097 1628 26153
rect 104 26067 130 26097
rect 1580 26067 1628 26097
rect 1618 26011 1628 26067
rect 104 25981 130 26011
rect 1580 25981 1628 26011
rect 1618 25925 1628 25981
rect 104 25895 130 25925
rect 1580 25895 1628 25925
rect 1618 25839 1628 25895
rect 104 25809 130 25839
rect 1580 25809 1628 25839
rect 1618 25753 1628 25809
rect 104 25723 130 25753
rect 1580 25723 1628 25753
rect 1618 25667 1628 25723
rect 104 25637 130 25667
rect 1580 25637 1628 25667
rect 1618 25581 1628 25637
rect 104 25551 130 25581
rect 1580 25551 1628 25581
rect 1618 25495 1628 25551
rect 104 25465 130 25495
rect 1580 25465 1628 25495
rect 1618 25409 1628 25465
rect 104 25379 130 25409
rect 1580 25379 1628 25409
rect 1618 25323 1628 25379
rect 104 25293 130 25323
rect 1580 25293 1628 25323
rect 1618 25237 1628 25293
rect 104 25207 130 25237
rect 1580 25207 1628 25237
rect 1618 25151 1628 25207
rect 104 25121 130 25151
rect 1580 25121 1628 25151
rect 1618 25065 1628 25121
rect 104 25035 130 25065
rect 1580 25035 1628 25065
rect 1618 24979 1628 25035
rect 104 24949 130 24979
rect 1580 24949 1628 24979
rect 1618 24893 1628 24949
rect 104 24863 130 24893
rect 1580 24863 1628 24893
rect 1618 24807 1628 24863
rect 104 24777 130 24807
rect 1580 24777 1628 24807
rect 1618 24721 1628 24777
rect 104 24691 130 24721
rect 1580 24691 1628 24721
rect 1618 24635 1628 24691
rect 104 24605 130 24635
rect 1580 24605 1628 24635
rect 1618 24549 1628 24605
rect 104 24519 130 24549
rect 1580 24519 1628 24549
rect 1618 24463 1628 24519
rect 104 24433 130 24463
rect 1580 24433 1628 24463
rect 1618 24377 1628 24433
rect 104 24347 130 24377
rect 1580 24347 1628 24377
rect 1618 24291 1628 24347
rect 104 24261 130 24291
rect 1580 24261 1628 24291
rect 1618 24205 1628 24261
rect 104 24175 130 24205
rect 1580 24175 1628 24205
rect 1618 24119 1628 24175
rect 104 24089 130 24119
rect 1580 24089 1628 24119
rect 1618 24033 1628 24089
rect 104 24003 130 24033
rect 1580 24003 1628 24033
rect 1618 23947 1628 24003
rect 104 23917 130 23947
rect 1580 23917 1628 23947
rect 1618 23861 1628 23917
rect 104 23831 130 23861
rect 1580 23831 1628 23861
rect 1618 23775 1628 23831
rect 104 23745 130 23775
rect 1580 23745 1628 23775
rect 1618 23689 1628 23745
rect 104 23659 130 23689
rect 1580 23659 1628 23689
rect 1618 23603 1628 23659
rect 104 23573 130 23603
rect 1580 23573 1628 23603
rect 1618 23517 1628 23573
rect 104 23487 130 23517
rect 1580 23487 1628 23517
rect 1618 23431 1628 23487
rect 104 23401 130 23431
rect 1580 23401 1628 23431
rect 1618 23345 1628 23401
rect 104 23315 130 23345
rect 1580 23315 1628 23345
rect 1618 23259 1628 23315
rect 104 23229 130 23259
rect 1580 23229 1628 23259
rect 1618 23173 1628 23229
rect 104 23143 130 23173
rect 1580 23143 1628 23173
rect 1618 23087 1628 23143
rect 104 23057 130 23087
rect 1580 23057 1628 23087
rect 1618 23001 1628 23057
rect 104 22971 130 23001
rect 1580 22971 1628 23001
rect 1618 22915 1628 22971
rect 104 22885 130 22915
rect 1580 22885 1628 22915
rect 1618 22829 1628 22885
rect 104 22799 130 22829
rect 1580 22799 1628 22829
rect 1618 22743 1628 22799
rect 104 22713 130 22743
rect 1580 22713 1628 22743
rect 1618 22657 1628 22713
rect 104 22627 130 22657
rect 1580 22627 1628 22657
rect 1618 22571 1628 22627
rect 104 22541 130 22571
rect 1580 22541 1628 22571
rect 1618 22485 1628 22541
rect 104 22455 130 22485
rect 1580 22455 1628 22485
rect 1618 22399 1628 22455
rect 104 22369 130 22399
rect 1580 22369 1628 22399
rect 1618 22313 1628 22369
rect 104 22283 130 22313
rect 1580 22283 1628 22313
rect 1618 22227 1628 22283
rect 104 22197 130 22227
rect 1580 22197 1628 22227
rect 1618 22141 1628 22197
rect 104 22111 130 22141
rect 1580 22111 1628 22141
rect 1618 22055 1628 22111
rect 104 22025 130 22055
rect 1580 22025 1628 22055
rect 1618 21969 1628 22025
rect 104 21939 130 21969
rect 1580 21939 1628 21969
rect 1618 21883 1628 21939
rect 104 21853 130 21883
rect 1580 21853 1628 21883
rect 1618 21797 1628 21853
rect 104 21767 130 21797
rect 1580 21767 1628 21797
rect 1618 21711 1628 21767
rect 104 21681 130 21711
rect 1580 21681 1628 21711
rect 1618 21625 1628 21681
rect 104 21595 130 21625
rect 1580 21595 1628 21625
rect 1618 21539 1628 21595
rect 104 21509 130 21539
rect 1580 21509 1628 21539
rect 1618 21453 1628 21509
rect 104 21423 130 21453
rect 1580 21423 1628 21453
rect 1618 21367 1628 21423
rect 104 21337 130 21367
rect 1580 21337 1628 21367
rect 1618 21281 1628 21337
rect 104 21251 130 21281
rect 1580 21251 1628 21281
rect 1618 21195 1628 21251
rect 104 21165 130 21195
rect 1580 21165 1628 21195
rect 1618 21109 1628 21165
rect 104 21079 130 21109
rect 1580 21079 1628 21109
rect 1618 21023 1628 21079
rect 104 20993 130 21023
rect 1580 20993 1628 21023
rect 1618 20937 1628 20993
rect 104 20907 130 20937
rect 1580 20907 1628 20937
rect 1618 20851 1628 20907
rect 104 20821 130 20851
rect 1580 20821 1628 20851
rect 1618 20765 1628 20821
rect 104 20735 130 20765
rect 1580 20735 1628 20765
rect 1618 20679 1628 20735
rect 104 20649 130 20679
rect 1580 20649 1628 20679
rect 1618 20593 1628 20649
rect 104 20563 130 20593
rect 1580 20563 1628 20593
rect 1618 20507 1628 20563
rect 104 20477 130 20507
rect 1580 20477 1628 20507
rect 1618 20421 1628 20477
rect 104 20391 130 20421
rect 1580 20391 1628 20421
rect 1618 20335 1628 20391
rect 104 20305 130 20335
rect 1580 20305 1628 20335
rect 1618 20249 1628 20305
rect 104 20219 130 20249
rect 1580 20219 1628 20249
rect 1618 20163 1628 20219
rect 104 20133 130 20163
rect 1580 20133 1628 20163
rect 1618 20077 1628 20133
rect 104 20047 130 20077
rect 1580 20047 1628 20077
rect 1618 19991 1628 20047
rect 104 19961 130 19991
rect 1580 19961 1628 19991
rect 1618 19905 1628 19961
rect 104 19875 130 19905
rect 1580 19875 1628 19905
rect 1618 19819 1628 19875
rect 104 19789 130 19819
rect 1580 19789 1628 19819
rect 1618 19733 1628 19789
rect 104 19703 130 19733
rect 1580 19703 1628 19733
rect 1618 19647 1628 19703
rect 104 19617 130 19647
rect 1580 19617 1628 19647
rect 1618 19561 1628 19617
rect 104 19531 130 19561
rect 1580 19531 1628 19561
rect 1618 19475 1628 19531
rect 104 19445 130 19475
rect 1580 19445 1628 19475
rect 1618 19389 1628 19445
rect 104 19359 130 19389
rect 1580 19359 1628 19389
rect 1618 19303 1628 19359
rect 104 19273 130 19303
rect 1580 19273 1628 19303
rect 1618 19217 1628 19273
rect 104 19187 130 19217
rect 1580 19187 1628 19217
rect 1618 19131 1628 19187
rect 104 19101 130 19131
rect 1580 19101 1628 19131
rect 1618 19045 1628 19101
rect 104 19015 130 19045
rect 1580 19015 1628 19045
rect 1618 18959 1628 19015
rect 104 18929 130 18959
rect 1580 18929 1628 18959
rect 1618 18873 1628 18929
rect 104 18843 130 18873
rect 1580 18843 1628 18873
rect 1618 18787 1628 18843
rect 104 18757 130 18787
rect 1580 18757 1628 18787
rect 1618 18701 1628 18757
rect 104 18671 130 18701
rect 1580 18671 1628 18701
rect 1618 18615 1628 18671
rect 104 18585 130 18615
rect 1580 18585 1628 18615
rect 1618 18529 1628 18585
rect 104 18499 130 18529
rect 1580 18499 1628 18529
rect 1618 18443 1628 18499
rect 104 18413 130 18443
rect 1580 18413 1628 18443
rect 1618 18357 1628 18413
rect 104 18327 130 18357
rect 1580 18327 1628 18357
rect 1618 18271 1628 18327
rect 104 18241 130 18271
rect 1580 18241 1628 18271
rect 1618 18185 1628 18241
rect 104 18155 130 18185
rect 1580 18155 1628 18185
rect 1618 18099 1628 18155
rect 104 18069 130 18099
rect 1580 18069 1628 18099
rect 1618 18013 1628 18069
rect 104 17983 130 18013
rect 1580 17983 1628 18013
rect 1618 17927 1628 17983
rect 104 17897 130 17927
rect 1580 17897 1628 17927
rect 1618 17841 1628 17897
rect 104 17811 130 17841
rect 1580 17811 1628 17841
rect 1618 17755 1628 17811
rect 104 17725 130 17755
rect 1580 17725 1628 17755
rect 1618 17669 1628 17725
rect 104 17639 130 17669
rect 1580 17639 1628 17669
rect 1618 17583 1628 17639
rect 104 17553 130 17583
rect 1580 17553 1628 17583
rect 1618 17497 1628 17553
rect 104 17467 130 17497
rect 1580 17467 1628 17497
rect 1618 17411 1628 17467
rect 104 17381 130 17411
rect 1580 17381 1628 17411
rect 1618 17325 1628 17381
rect 104 17295 130 17325
rect 1580 17295 1628 17325
rect 1618 17239 1628 17295
rect 104 17209 130 17239
rect 1580 17209 1628 17239
rect 1618 17153 1628 17209
rect 104 17123 130 17153
rect 1580 17123 1628 17153
rect 1618 17067 1628 17123
rect 104 17037 130 17067
rect 1580 17037 1628 17067
rect 1618 16981 1628 17037
rect 104 16951 130 16981
rect 1580 16951 1628 16981
rect 1618 16895 1628 16951
rect 104 16865 130 16895
rect 1580 16865 1628 16895
rect 1618 16809 1628 16865
rect 104 16779 130 16809
rect 1580 16779 1628 16809
rect 1618 16723 1628 16779
rect 104 16693 130 16723
rect 1580 16693 1628 16723
rect 1618 16637 1628 16693
rect 104 16607 130 16637
rect 1580 16607 1628 16637
rect 1618 16551 1628 16607
rect 104 16521 130 16551
rect 1580 16521 1628 16551
rect 1618 16465 1628 16521
rect 104 16435 130 16465
rect 1580 16435 1628 16465
rect 1618 16379 1628 16435
rect 104 16349 130 16379
rect 1580 16349 1628 16379
rect 1618 16293 1628 16349
rect 104 16263 130 16293
rect 1580 16263 1628 16293
rect 1618 16207 1628 16263
rect 104 16177 130 16207
rect 1580 16177 1628 16207
rect 1618 16121 1628 16177
rect 104 16091 130 16121
rect 1580 16091 1628 16121
rect 1618 16035 1628 16091
rect 104 16005 130 16035
rect 1580 16005 1628 16035
rect 1618 15949 1628 16005
rect 104 15919 130 15949
rect 1580 15919 1628 15949
rect 1618 15863 1628 15919
rect 104 15833 130 15863
rect 1580 15833 1628 15863
rect 1618 15777 1628 15833
rect 104 15747 130 15777
rect 1580 15747 1628 15777
rect 1618 15691 1628 15747
rect 104 15661 130 15691
rect 1580 15661 1628 15691
rect 1618 15605 1628 15661
rect 104 15575 130 15605
rect 1580 15575 1628 15605
rect 1618 15519 1628 15575
rect 104 15489 130 15519
rect 1580 15489 1628 15519
rect 1618 15433 1628 15489
rect 104 15403 130 15433
rect 1580 15403 1628 15433
rect 1618 15347 1628 15403
rect 104 15317 130 15347
rect 1580 15317 1628 15347
rect 1618 15261 1628 15317
rect 104 15231 130 15261
rect 1580 15231 1628 15261
rect 1618 15175 1628 15231
rect 104 15145 130 15175
rect 1580 15145 1628 15175
rect 1618 15089 1628 15145
rect 104 15059 130 15089
rect 1580 15059 1628 15089
rect 1618 15003 1628 15059
rect 104 14973 130 15003
rect 1580 14973 1628 15003
rect 1618 14917 1628 14973
rect 104 14887 130 14917
rect 1580 14887 1628 14917
rect 1618 14831 1628 14887
rect 104 14801 130 14831
rect 1580 14801 1628 14831
rect 1618 14745 1628 14801
rect 104 14715 130 14745
rect 1580 14715 1628 14745
rect 1618 14659 1628 14715
rect 104 14629 130 14659
rect 1580 14629 1628 14659
rect 1618 14573 1628 14629
rect 104 14543 130 14573
rect 1580 14543 1628 14573
rect 1618 14487 1628 14543
rect 104 14457 130 14487
rect 1580 14457 1628 14487
rect 1618 14401 1628 14457
rect 104 14371 130 14401
rect 1580 14371 1628 14401
rect 1618 14315 1628 14371
rect 104 14285 130 14315
rect 1580 14285 1628 14315
rect 1618 14229 1628 14285
rect 104 14199 130 14229
rect 1580 14199 1628 14229
rect 1618 14143 1628 14199
rect 104 14113 130 14143
rect 1580 14113 1628 14143
rect 1618 14057 1628 14113
rect 104 14027 130 14057
rect 1580 14027 1628 14057
rect 1618 13971 1628 14027
rect 104 13941 130 13971
rect 1580 13941 1628 13971
rect 1618 13885 1628 13941
rect 104 13855 130 13885
rect 1580 13855 1628 13885
rect 1618 13799 1628 13855
rect 104 13769 130 13799
rect 1580 13769 1628 13799
rect 1618 13713 1628 13769
rect 104 13683 130 13713
rect 1580 13683 1628 13713
rect 1618 13627 1628 13683
rect 104 13597 130 13627
rect 1580 13597 1628 13627
rect 1618 13541 1628 13597
rect 104 13511 130 13541
rect 1580 13511 1628 13541
rect 1618 13455 1628 13511
rect 104 13425 130 13455
rect 1580 13425 1628 13455
rect 1618 13369 1628 13425
rect 104 13339 130 13369
rect 1580 13339 1628 13369
rect 1618 13283 1628 13339
rect 104 13253 130 13283
rect 1580 13253 1628 13283
rect 1618 13197 1628 13253
rect 104 13167 130 13197
rect 1580 13167 1628 13197
rect 1618 13111 1628 13167
rect 104 13081 130 13111
rect 1580 13081 1628 13111
rect 1618 13025 1628 13081
rect 104 12995 130 13025
rect 1580 12995 1628 13025
rect 1618 12939 1628 12995
rect 104 12909 130 12939
rect 1580 12909 1628 12939
rect 1618 12853 1628 12909
rect 104 12823 130 12853
rect 1580 12823 1628 12853
rect 1618 12767 1628 12823
rect 104 12737 130 12767
rect 1580 12737 1628 12767
rect 1618 12681 1628 12737
rect 104 12651 130 12681
rect 1580 12651 1628 12681
rect 1618 12595 1628 12651
rect 104 12565 130 12595
rect 1580 12565 1628 12595
rect 1618 12509 1628 12565
rect 104 12479 130 12509
rect 1580 12479 1628 12509
rect 1618 12423 1628 12479
rect 104 12393 130 12423
rect 1580 12393 1628 12423
rect 1618 12337 1628 12393
rect 104 12307 130 12337
rect 1580 12307 1628 12337
rect 1618 12251 1628 12307
rect 104 12221 130 12251
rect 1580 12221 1628 12251
rect 1618 12165 1628 12221
rect 104 12135 130 12165
rect 1580 12135 1628 12165
rect 1618 12079 1628 12135
rect 104 12049 130 12079
rect 1580 12049 1628 12079
rect 1618 11993 1628 12049
rect 104 11963 130 11993
rect 1580 11963 1628 11993
rect 1618 11907 1628 11963
rect 104 11877 130 11907
rect 1580 11877 1628 11907
rect 1618 11821 1628 11877
rect 104 11791 130 11821
rect 1580 11791 1628 11821
rect 1618 11735 1628 11791
rect 104 11705 130 11735
rect 1580 11705 1628 11735
rect 1618 11649 1628 11705
rect 104 11619 130 11649
rect 1580 11619 1628 11649
rect 1618 11563 1628 11619
rect 104 11533 130 11563
rect 1580 11533 1628 11563
rect 1618 11477 1628 11533
rect 104 11447 130 11477
rect 1580 11447 1628 11477
rect 1618 11391 1628 11447
rect 104 11361 130 11391
rect 1580 11361 1628 11391
rect 1618 11305 1628 11361
rect 104 11275 130 11305
rect 1580 11275 1628 11305
rect 1618 11219 1628 11275
rect 104 11189 130 11219
rect 1580 11189 1628 11219
rect 1618 11133 1628 11189
rect 104 11103 130 11133
rect 1580 11103 1628 11133
rect 1618 11047 1628 11103
rect 104 11017 130 11047
rect 1580 11017 1628 11047
rect 1618 10961 1628 11017
rect 104 10931 130 10961
rect 1580 10931 1628 10961
rect 1618 10875 1628 10931
rect 104 10845 130 10875
rect 1580 10845 1628 10875
rect 1618 10789 1628 10845
rect 104 10759 130 10789
rect 1580 10759 1628 10789
rect 1618 10703 1628 10759
rect 104 10673 130 10703
rect 1580 10673 1628 10703
rect 1618 10617 1628 10673
rect 104 10587 130 10617
rect 1580 10587 1628 10617
rect 1618 10531 1628 10587
rect 104 10501 130 10531
rect 1580 10501 1628 10531
rect 1618 10445 1628 10501
rect 104 10415 130 10445
rect 1580 10415 1628 10445
rect 1618 10359 1628 10415
rect 104 10329 130 10359
rect 1580 10329 1628 10359
rect 1618 10273 1628 10329
rect 104 10243 130 10273
rect 1580 10243 1628 10273
rect 1618 10187 1628 10243
rect 104 10157 130 10187
rect 1580 10157 1628 10187
rect 1618 10101 1628 10157
rect 104 10071 130 10101
rect 1580 10071 1628 10101
rect 1618 10015 1628 10071
rect 104 9985 130 10015
rect 1580 9985 1628 10015
rect 1618 9929 1628 9985
rect 104 9899 130 9929
rect 1580 9899 1628 9929
rect 1618 9843 1628 9899
rect 104 9813 130 9843
rect 1580 9813 1628 9843
rect 1618 9757 1628 9813
rect 104 9727 130 9757
rect 1580 9727 1628 9757
rect 1618 9671 1628 9727
rect 104 9641 130 9671
rect 1580 9641 1628 9671
rect 1618 9585 1628 9641
rect 104 9555 130 9585
rect 1580 9555 1628 9585
rect 1618 9499 1628 9555
rect 104 9469 130 9499
rect 1580 9469 1628 9499
rect 1618 9413 1628 9469
rect 104 9383 130 9413
rect 1580 9383 1628 9413
rect 1618 9327 1628 9383
rect 104 9297 130 9327
rect 1580 9297 1628 9327
rect 1618 9241 1628 9297
rect 104 9211 130 9241
rect 1580 9211 1628 9241
rect 1618 9155 1628 9211
rect 104 9125 130 9155
rect 1580 9125 1628 9155
rect 1618 9069 1628 9125
rect 104 9039 130 9069
rect 1580 9039 1628 9069
rect 1618 8983 1628 9039
rect 104 8953 130 8983
rect 1580 8953 1628 8983
rect 1618 8897 1628 8953
rect 104 8867 130 8897
rect 1580 8867 1628 8897
rect 1618 8811 1628 8867
rect 104 8781 130 8811
rect 1580 8781 1628 8811
rect 1618 8725 1628 8781
rect 104 8695 130 8725
rect 1580 8695 1628 8725
rect 1618 8639 1628 8695
rect 104 8609 130 8639
rect 1580 8609 1628 8639
rect 1618 8553 1628 8609
rect 104 8523 130 8553
rect 1580 8523 1628 8553
rect 1618 8467 1628 8523
rect 104 8437 130 8467
rect 1580 8437 1628 8467
rect 1618 8381 1628 8437
rect 104 8351 130 8381
rect 1580 8351 1628 8381
rect 1618 8295 1628 8351
rect 104 8265 130 8295
rect 1580 8265 1628 8295
rect 1618 8209 1628 8265
rect 104 8179 130 8209
rect 1580 8179 1628 8209
rect 1618 8123 1628 8179
rect 104 8093 130 8123
rect 1580 8093 1628 8123
rect 1618 8037 1628 8093
rect 104 8007 130 8037
rect 1580 8007 1628 8037
rect 1618 7951 1628 8007
rect 104 7921 130 7951
rect 1580 7921 1628 7951
rect 1618 7865 1628 7921
rect 104 7835 130 7865
rect 1580 7835 1628 7865
rect 1618 7779 1628 7835
rect 104 7749 130 7779
rect 1580 7749 1628 7779
rect 1618 7693 1628 7749
rect 104 7663 130 7693
rect 1580 7663 1628 7693
rect 1618 7607 1628 7663
rect 104 7577 130 7607
rect 1580 7577 1628 7607
rect 1618 7521 1628 7577
rect 104 7491 130 7521
rect 1580 7491 1628 7521
rect 1618 7435 1628 7491
rect 104 7405 130 7435
rect 1580 7405 1628 7435
rect 1618 7349 1628 7405
rect 104 7319 130 7349
rect 1580 7319 1628 7349
rect 1618 7263 1628 7319
rect 104 7233 130 7263
rect 1580 7233 1628 7263
rect 1618 7177 1628 7233
rect 104 7147 130 7177
rect 1580 7147 1628 7177
rect 1618 7091 1628 7147
rect 104 7061 130 7091
rect 1580 7061 1628 7091
rect 1618 7005 1628 7061
rect 104 6975 130 7005
rect 1580 6975 1628 7005
rect 1618 6919 1628 6975
rect 104 6889 130 6919
rect 1580 6889 1628 6919
rect 1618 6833 1628 6889
rect 104 6803 130 6833
rect 1580 6803 1628 6833
rect 1618 6747 1628 6803
rect 104 6717 130 6747
rect 1580 6717 1628 6747
rect 1618 6661 1628 6717
rect 104 6631 130 6661
rect 1580 6631 1628 6661
rect 1618 6575 1628 6631
rect 104 6545 130 6575
rect 1580 6545 1628 6575
rect 1618 6489 1628 6545
rect 104 6459 130 6489
rect 1580 6459 1628 6489
rect 1618 6403 1628 6459
rect 104 6373 130 6403
rect 1580 6373 1628 6403
rect 1618 6317 1628 6373
rect 104 6287 130 6317
rect 1580 6287 1628 6317
rect 1618 6231 1628 6287
rect 104 6201 130 6231
rect 1580 6201 1628 6231
rect 1618 6145 1628 6201
rect 104 6115 130 6145
rect 1580 6115 1628 6145
rect 1618 6059 1628 6115
rect 104 6029 130 6059
rect 1580 6029 1628 6059
rect 1618 5973 1628 6029
rect 104 5943 130 5973
rect 1580 5943 1628 5973
rect 1618 5887 1628 5943
rect 104 5857 130 5887
rect 1580 5857 1628 5887
rect 1618 5801 1628 5857
rect 104 5771 130 5801
rect 1580 5771 1628 5801
rect 1618 5715 1628 5771
rect 104 5685 130 5715
rect 1580 5685 1628 5715
rect 1618 5629 1628 5685
rect 104 5599 130 5629
rect 1580 5599 1628 5629
rect 1618 5543 1628 5599
rect 104 5513 130 5543
rect 1580 5513 1628 5543
rect 1618 5457 1628 5513
rect 104 5427 130 5457
rect 1580 5427 1628 5457
rect 1618 5371 1628 5427
rect 104 5341 130 5371
rect 1580 5341 1628 5371
rect 1618 5285 1628 5341
rect 104 5255 130 5285
rect 1580 5255 1628 5285
rect 1618 5199 1628 5255
rect 104 5169 130 5199
rect 1580 5169 1628 5199
rect 1618 5113 1628 5169
rect 104 5083 130 5113
rect 1580 5083 1628 5113
rect 1618 5027 1628 5083
rect 104 4997 130 5027
rect 1580 4997 1628 5027
rect 1618 4941 1628 4997
rect 104 4911 130 4941
rect 1580 4911 1628 4941
rect 1618 4855 1628 4911
rect 104 4825 130 4855
rect 1580 4825 1628 4855
rect 1618 4769 1628 4825
rect 104 4739 130 4769
rect 1580 4739 1628 4769
rect 1618 4683 1628 4739
rect 104 4653 130 4683
rect 1580 4653 1628 4683
rect 1618 4597 1628 4653
rect 104 4567 130 4597
rect 1580 4567 1628 4597
rect 1618 4511 1628 4567
rect 104 4481 130 4511
rect 1580 4481 1628 4511
rect 1618 4425 1628 4481
rect 104 4395 130 4425
rect 1580 4395 1628 4425
rect 1618 4339 1628 4395
rect 104 4309 130 4339
rect 1580 4309 1628 4339
rect 1618 4253 1628 4309
rect 104 4223 130 4253
rect 1580 4223 1628 4253
rect 1618 4167 1628 4223
rect 104 4137 130 4167
rect 1580 4137 1628 4167
rect 1618 4081 1628 4137
rect 104 4051 130 4081
rect 1580 4051 1628 4081
rect 1618 3995 1628 4051
rect 104 3965 130 3995
rect 1580 3965 1628 3995
rect 1618 3909 1628 3965
rect 104 3879 130 3909
rect 1580 3879 1628 3909
rect 1618 3823 1628 3879
rect 104 3793 130 3823
rect 1580 3793 1628 3823
rect 1618 3737 1628 3793
rect 104 3707 130 3737
rect 1580 3707 1628 3737
rect 1618 3651 1628 3707
rect 104 3621 130 3651
rect 1580 3621 1628 3651
rect 1618 3565 1628 3621
rect 104 3535 130 3565
rect 1580 3535 1628 3565
rect 1618 3479 1628 3535
rect 104 3449 130 3479
rect 1580 3449 1628 3479
rect 1618 3393 1628 3449
rect 104 3363 130 3393
rect 1580 3363 1628 3393
rect 1618 3307 1628 3363
rect 104 3277 130 3307
rect 1580 3277 1628 3307
rect 1618 3221 1628 3277
rect 104 3191 130 3221
rect 1580 3191 1628 3221
rect 1618 3135 1628 3191
rect 104 3105 130 3135
rect 1580 3105 1628 3135
rect 1618 3049 1628 3105
rect 104 3019 130 3049
rect 1580 3019 1628 3049
rect 1618 2963 1628 3019
rect 104 2933 130 2963
rect 1580 2933 1628 2963
rect 1618 2877 1628 2933
rect 104 2847 130 2877
rect 1580 2847 1628 2877
rect 1618 2791 1628 2847
rect 104 2761 130 2791
rect 1580 2761 1628 2791
rect 1618 2705 1628 2761
rect 104 2675 130 2705
rect 1580 2675 1628 2705
rect 1618 2619 1628 2675
rect 104 2589 130 2619
rect 1580 2589 1628 2619
rect 1618 2533 1628 2589
rect 104 2503 130 2533
rect 1580 2503 1628 2533
rect 1618 2447 1628 2503
rect 104 2417 130 2447
rect 1580 2417 1628 2447
rect 1618 2361 1628 2417
rect 104 2331 130 2361
rect 1580 2331 1628 2361
rect 1618 2275 1628 2331
rect 104 2245 130 2275
rect 1580 2245 1628 2275
rect 1618 2189 1628 2245
rect 104 2159 130 2189
rect 1580 2159 1628 2189
rect 1618 2103 1628 2159
rect 104 2073 130 2103
rect 1580 2073 1628 2103
rect 1618 2017 1628 2073
rect 104 1987 130 2017
rect 1580 1987 1628 2017
rect 1618 1931 1628 1987
rect 104 1901 130 1931
rect 1580 1901 1628 1931
rect 1618 1845 1628 1901
rect 104 1815 130 1845
rect 1580 1815 1628 1845
rect 1618 1759 1628 1815
rect 104 1729 130 1759
rect 1580 1729 1628 1759
rect 1618 1673 1628 1729
rect 104 1643 130 1673
rect 1580 1643 1628 1673
rect 1618 1587 1628 1643
rect 104 1557 130 1587
rect 1580 1557 1628 1587
rect 1618 1501 1628 1557
rect 104 1471 130 1501
rect 1580 1471 1628 1501
rect 1618 1415 1628 1471
rect 104 1385 130 1415
rect 1580 1385 1628 1415
rect 1618 1329 1628 1385
rect 104 1299 130 1329
rect 1580 1299 1628 1329
rect 1618 1243 1628 1299
rect 104 1213 130 1243
rect 1580 1213 1628 1243
rect 1618 1157 1628 1213
rect 104 1127 130 1157
rect 1580 1127 1628 1157
rect 1618 1071 1628 1127
rect 104 1041 130 1071
rect 1580 1041 1628 1071
rect 1618 985 1628 1041
rect 104 955 130 985
rect 1580 955 1628 985
rect 1618 899 1628 955
rect 104 869 130 899
rect 1580 869 1628 899
rect 1618 813 1628 869
rect 104 783 130 813
rect 1580 783 1628 813
rect 1618 727 1628 783
rect 104 697 130 727
rect 1580 697 1628 727
rect 1618 641 1628 697
rect 104 611 130 641
rect 1580 611 1628 641
rect 1618 555 1628 611
rect 104 525 130 555
rect 1580 525 1628 555
rect 1618 469 1628 525
rect 104 439 130 469
rect 1580 439 1628 469
rect 1618 383 1628 439
rect 104 353 130 383
rect 1580 353 1628 383
rect 1618 297 1628 353
rect 104 267 130 297
rect 1580 267 1628 297
rect 1618 211 1628 267
rect 104 181 130 211
rect 1580 181 1628 211
rect 1618 179 1628 181
rect 1662 179 1672 100059
rect 1618 163 1672 179
<< polycont >>
rect 1628 179 1662 100059
<< locali >>
rect 36 100168 100 100202
rect 1680 100168 1744 100202
rect 36 100138 70 100168
rect 1710 100138 1744 100168
rect 122 100068 138 100102
rect 1572 100068 1588 100102
rect 1628 100059 1662 100075
rect 122 99982 138 100016
rect 1572 99982 1588 100016
rect 122 99896 138 99930
rect 1572 99896 1588 99930
rect 122 99810 138 99844
rect 1572 99810 1588 99844
rect 122 99724 138 99758
rect 1572 99724 1588 99758
rect 122 99638 138 99672
rect 1572 99638 1588 99672
rect 122 99552 138 99586
rect 1572 99552 1588 99586
rect 122 99466 138 99500
rect 1572 99466 1588 99500
rect 122 99380 138 99414
rect 1572 99380 1588 99414
rect 122 99294 138 99328
rect 1572 99294 1588 99328
rect 122 99208 138 99242
rect 1572 99208 1588 99242
rect 122 99122 138 99156
rect 1572 99122 1588 99156
rect 122 99036 138 99070
rect 1572 99036 1588 99070
rect 122 98950 138 98984
rect 1572 98950 1588 98984
rect 122 98864 138 98898
rect 1572 98864 1588 98898
rect 122 98778 138 98812
rect 1572 98778 1588 98812
rect 122 98692 138 98726
rect 1572 98692 1588 98726
rect 122 98606 138 98640
rect 1572 98606 1588 98640
rect 122 98520 138 98554
rect 1572 98520 1588 98554
rect 122 98434 138 98468
rect 1572 98434 1588 98468
rect 122 98348 138 98382
rect 1572 98348 1588 98382
rect 122 98262 138 98296
rect 1572 98262 1588 98296
rect 122 98176 138 98210
rect 1572 98176 1588 98210
rect 122 98090 138 98124
rect 1572 98090 1588 98124
rect 122 98004 138 98038
rect 1572 98004 1588 98038
rect 122 97918 138 97952
rect 1572 97918 1588 97952
rect 122 97832 138 97866
rect 1572 97832 1588 97866
rect 122 97746 138 97780
rect 1572 97746 1588 97780
rect 122 97660 138 97694
rect 1572 97660 1588 97694
rect 122 97574 138 97608
rect 1572 97574 1588 97608
rect 122 97488 138 97522
rect 1572 97488 1588 97522
rect 122 97402 138 97436
rect 1572 97402 1588 97436
rect 122 97316 138 97350
rect 1572 97316 1588 97350
rect 122 97230 138 97264
rect 1572 97230 1588 97264
rect 122 97144 138 97178
rect 1572 97144 1588 97178
rect 122 97058 138 97092
rect 1572 97058 1588 97092
rect 122 96972 138 97006
rect 1572 96972 1588 97006
rect 122 96886 138 96920
rect 1572 96886 1588 96920
rect 122 96800 138 96834
rect 1572 96800 1588 96834
rect 122 96714 138 96748
rect 1572 96714 1588 96748
rect 122 96628 138 96662
rect 1572 96628 1588 96662
rect 122 96542 138 96576
rect 1572 96542 1588 96576
rect 122 96456 138 96490
rect 1572 96456 1588 96490
rect 122 96370 138 96404
rect 1572 96370 1588 96404
rect 122 96284 138 96318
rect 1572 96284 1588 96318
rect 122 96198 138 96232
rect 1572 96198 1588 96232
rect 122 96112 138 96146
rect 1572 96112 1588 96146
rect 122 96026 138 96060
rect 1572 96026 1588 96060
rect 122 95940 138 95974
rect 1572 95940 1588 95974
rect 122 95854 138 95888
rect 1572 95854 1588 95888
rect 122 95768 138 95802
rect 1572 95768 1588 95802
rect 122 95682 138 95716
rect 1572 95682 1588 95716
rect 122 95596 138 95630
rect 1572 95596 1588 95630
rect 122 95510 138 95544
rect 1572 95510 1588 95544
rect 122 95424 138 95458
rect 1572 95424 1588 95458
rect 122 95338 138 95372
rect 1572 95338 1588 95372
rect 122 95252 138 95286
rect 1572 95252 1588 95286
rect 122 95166 138 95200
rect 1572 95166 1588 95200
rect 122 95080 138 95114
rect 1572 95080 1588 95114
rect 122 94994 138 95028
rect 1572 94994 1588 95028
rect 122 94908 138 94942
rect 1572 94908 1588 94942
rect 122 94822 138 94856
rect 1572 94822 1588 94856
rect 122 94736 138 94770
rect 1572 94736 1588 94770
rect 122 94650 138 94684
rect 1572 94650 1588 94684
rect 122 94564 138 94598
rect 1572 94564 1588 94598
rect 122 94478 138 94512
rect 1572 94478 1588 94512
rect 122 94392 138 94426
rect 1572 94392 1588 94426
rect 122 94306 138 94340
rect 1572 94306 1588 94340
rect 122 94220 138 94254
rect 1572 94220 1588 94254
rect 122 94134 138 94168
rect 1572 94134 1588 94168
rect 122 94048 138 94082
rect 1572 94048 1588 94082
rect 122 93962 138 93996
rect 1572 93962 1588 93996
rect 122 93876 138 93910
rect 1572 93876 1588 93910
rect 122 93790 138 93824
rect 1572 93790 1588 93824
rect 122 93704 138 93738
rect 1572 93704 1588 93738
rect 122 93618 138 93652
rect 1572 93618 1588 93652
rect 122 93532 138 93566
rect 1572 93532 1588 93566
rect 122 93446 138 93480
rect 1572 93446 1588 93480
rect 122 93360 138 93394
rect 1572 93360 1588 93394
rect 122 93274 138 93308
rect 1572 93274 1588 93308
rect 122 93188 138 93222
rect 1572 93188 1588 93222
rect 122 93102 138 93136
rect 1572 93102 1588 93136
rect 122 93016 138 93050
rect 1572 93016 1588 93050
rect 122 92930 138 92964
rect 1572 92930 1588 92964
rect 122 92844 138 92878
rect 1572 92844 1588 92878
rect 122 92758 138 92792
rect 1572 92758 1588 92792
rect 122 92672 138 92706
rect 1572 92672 1588 92706
rect 122 92586 138 92620
rect 1572 92586 1588 92620
rect 122 92500 138 92534
rect 1572 92500 1588 92534
rect 122 92414 138 92448
rect 1572 92414 1588 92448
rect 122 92328 138 92362
rect 1572 92328 1588 92362
rect 122 92242 138 92276
rect 1572 92242 1588 92276
rect 122 92156 138 92190
rect 1572 92156 1588 92190
rect 122 92070 138 92104
rect 1572 92070 1588 92104
rect 122 91984 138 92018
rect 1572 91984 1588 92018
rect 122 91898 138 91932
rect 1572 91898 1588 91932
rect 122 91812 138 91846
rect 1572 91812 1588 91846
rect 122 91726 138 91760
rect 1572 91726 1588 91760
rect 122 91640 138 91674
rect 1572 91640 1588 91674
rect 122 91554 138 91588
rect 1572 91554 1588 91588
rect 122 91468 138 91502
rect 1572 91468 1588 91502
rect 122 91382 138 91416
rect 1572 91382 1588 91416
rect 122 91296 138 91330
rect 1572 91296 1588 91330
rect 122 91210 138 91244
rect 1572 91210 1588 91244
rect 122 91124 138 91158
rect 1572 91124 1588 91158
rect 122 91038 138 91072
rect 1572 91038 1588 91072
rect 122 90952 138 90986
rect 1572 90952 1588 90986
rect 122 90866 138 90900
rect 1572 90866 1588 90900
rect 122 90780 138 90814
rect 1572 90780 1588 90814
rect 122 90694 138 90728
rect 1572 90694 1588 90728
rect 122 90608 138 90642
rect 1572 90608 1588 90642
rect 122 90522 138 90556
rect 1572 90522 1588 90556
rect 122 90436 138 90470
rect 1572 90436 1588 90470
rect 122 90350 138 90384
rect 1572 90350 1588 90384
rect 122 90264 138 90298
rect 1572 90264 1588 90298
rect 122 90178 138 90212
rect 1572 90178 1588 90212
rect 122 90092 138 90126
rect 1572 90092 1588 90126
rect 122 90006 138 90040
rect 1572 90006 1588 90040
rect 122 89920 138 89954
rect 1572 89920 1588 89954
rect 122 89834 138 89868
rect 1572 89834 1588 89868
rect 122 89748 138 89782
rect 1572 89748 1588 89782
rect 122 89662 138 89696
rect 1572 89662 1588 89696
rect 122 89576 138 89610
rect 1572 89576 1588 89610
rect 122 89490 138 89524
rect 1572 89490 1588 89524
rect 122 89404 138 89438
rect 1572 89404 1588 89438
rect 122 89318 138 89352
rect 1572 89318 1588 89352
rect 122 89232 138 89266
rect 1572 89232 1588 89266
rect 122 89146 138 89180
rect 1572 89146 1588 89180
rect 122 89060 138 89094
rect 1572 89060 1588 89094
rect 122 88974 138 89008
rect 1572 88974 1588 89008
rect 122 88888 138 88922
rect 1572 88888 1588 88922
rect 122 88802 138 88836
rect 1572 88802 1588 88836
rect 122 88716 138 88750
rect 1572 88716 1588 88750
rect 122 88630 138 88664
rect 1572 88630 1588 88664
rect 122 88544 138 88578
rect 1572 88544 1588 88578
rect 122 88458 138 88492
rect 1572 88458 1588 88492
rect 122 88372 138 88406
rect 1572 88372 1588 88406
rect 122 88286 138 88320
rect 1572 88286 1588 88320
rect 122 88200 138 88234
rect 1572 88200 1588 88234
rect 122 88114 138 88148
rect 1572 88114 1588 88148
rect 122 88028 138 88062
rect 1572 88028 1588 88062
rect 122 87942 138 87976
rect 1572 87942 1588 87976
rect 122 87856 138 87890
rect 1572 87856 1588 87890
rect 122 87770 138 87804
rect 1572 87770 1588 87804
rect 122 87684 138 87718
rect 1572 87684 1588 87718
rect 122 87598 138 87632
rect 1572 87598 1588 87632
rect 122 87512 138 87546
rect 1572 87512 1588 87546
rect 122 87426 138 87460
rect 1572 87426 1588 87460
rect 122 87340 138 87374
rect 1572 87340 1588 87374
rect 122 87254 138 87288
rect 1572 87254 1588 87288
rect 122 87168 138 87202
rect 1572 87168 1588 87202
rect 122 87082 138 87116
rect 1572 87082 1588 87116
rect 122 86996 138 87030
rect 1572 86996 1588 87030
rect 122 86910 138 86944
rect 1572 86910 1588 86944
rect 122 86824 138 86858
rect 1572 86824 1588 86858
rect 122 86738 138 86772
rect 1572 86738 1588 86772
rect 122 86652 138 86686
rect 1572 86652 1588 86686
rect 122 86566 138 86600
rect 1572 86566 1588 86600
rect 122 86480 138 86514
rect 1572 86480 1588 86514
rect 122 86394 138 86428
rect 1572 86394 1588 86428
rect 122 86308 138 86342
rect 1572 86308 1588 86342
rect 122 86222 138 86256
rect 1572 86222 1588 86256
rect 122 86136 138 86170
rect 1572 86136 1588 86170
rect 122 86050 138 86084
rect 1572 86050 1588 86084
rect 122 85964 138 85998
rect 1572 85964 1588 85998
rect 122 85878 138 85912
rect 1572 85878 1588 85912
rect 122 85792 138 85826
rect 1572 85792 1588 85826
rect 122 85706 138 85740
rect 1572 85706 1588 85740
rect 122 85620 138 85654
rect 1572 85620 1588 85654
rect 122 85534 138 85568
rect 1572 85534 1588 85568
rect 122 85448 138 85482
rect 1572 85448 1588 85482
rect 122 85362 138 85396
rect 1572 85362 1588 85396
rect 122 85276 138 85310
rect 1572 85276 1588 85310
rect 122 85190 138 85224
rect 1572 85190 1588 85224
rect 122 85104 138 85138
rect 1572 85104 1588 85138
rect 122 85018 138 85052
rect 1572 85018 1588 85052
rect 122 84932 138 84966
rect 1572 84932 1588 84966
rect 122 84846 138 84880
rect 1572 84846 1588 84880
rect 122 84760 138 84794
rect 1572 84760 1588 84794
rect 122 84674 138 84708
rect 1572 84674 1588 84708
rect 122 84588 138 84622
rect 1572 84588 1588 84622
rect 122 84502 138 84536
rect 1572 84502 1588 84536
rect 122 84416 138 84450
rect 1572 84416 1588 84450
rect 122 84330 138 84364
rect 1572 84330 1588 84364
rect 122 84244 138 84278
rect 1572 84244 1588 84278
rect 122 84158 138 84192
rect 1572 84158 1588 84192
rect 122 84072 138 84106
rect 1572 84072 1588 84106
rect 122 83986 138 84020
rect 1572 83986 1588 84020
rect 122 83900 138 83934
rect 1572 83900 1588 83934
rect 122 83814 138 83848
rect 1572 83814 1588 83848
rect 122 83728 138 83762
rect 1572 83728 1588 83762
rect 122 83642 138 83676
rect 1572 83642 1588 83676
rect 122 83556 138 83590
rect 1572 83556 1588 83590
rect 122 83470 138 83504
rect 1572 83470 1588 83504
rect 122 83384 138 83418
rect 1572 83384 1588 83418
rect 122 83298 138 83332
rect 1572 83298 1588 83332
rect 122 83212 138 83246
rect 1572 83212 1588 83246
rect 122 83126 138 83160
rect 1572 83126 1588 83160
rect 122 83040 138 83074
rect 1572 83040 1588 83074
rect 122 82954 138 82988
rect 1572 82954 1588 82988
rect 122 82868 138 82902
rect 1572 82868 1588 82902
rect 122 82782 138 82816
rect 1572 82782 1588 82816
rect 122 82696 138 82730
rect 1572 82696 1588 82730
rect 122 82610 138 82644
rect 1572 82610 1588 82644
rect 122 82524 138 82558
rect 1572 82524 1588 82558
rect 122 82438 138 82472
rect 1572 82438 1588 82472
rect 122 82352 138 82386
rect 1572 82352 1588 82386
rect 122 82266 138 82300
rect 1572 82266 1588 82300
rect 122 82180 138 82214
rect 1572 82180 1588 82214
rect 122 82094 138 82128
rect 1572 82094 1588 82128
rect 122 82008 138 82042
rect 1572 82008 1588 82042
rect 122 81922 138 81956
rect 1572 81922 1588 81956
rect 122 81836 138 81870
rect 1572 81836 1588 81870
rect 122 81750 138 81784
rect 1572 81750 1588 81784
rect 122 81664 138 81698
rect 1572 81664 1588 81698
rect 122 81578 138 81612
rect 1572 81578 1588 81612
rect 122 81492 138 81526
rect 1572 81492 1588 81526
rect 122 81406 138 81440
rect 1572 81406 1588 81440
rect 122 81320 138 81354
rect 1572 81320 1588 81354
rect 122 81234 138 81268
rect 1572 81234 1588 81268
rect 122 81148 138 81182
rect 1572 81148 1588 81182
rect 122 81062 138 81096
rect 1572 81062 1588 81096
rect 122 80976 138 81010
rect 1572 80976 1588 81010
rect 122 80890 138 80924
rect 1572 80890 1588 80924
rect 122 80804 138 80838
rect 1572 80804 1588 80838
rect 122 80718 138 80752
rect 1572 80718 1588 80752
rect 122 80632 138 80666
rect 1572 80632 1588 80666
rect 122 80546 138 80580
rect 1572 80546 1588 80580
rect 122 80460 138 80494
rect 1572 80460 1588 80494
rect 122 80374 138 80408
rect 1572 80374 1588 80408
rect 122 80288 138 80322
rect 1572 80288 1588 80322
rect 122 80202 138 80236
rect 1572 80202 1588 80236
rect 122 80116 138 80150
rect 1572 80116 1588 80150
rect 122 80030 138 80064
rect 1572 80030 1588 80064
rect 122 79944 138 79978
rect 1572 79944 1588 79978
rect 122 79858 138 79892
rect 1572 79858 1588 79892
rect 122 79772 138 79806
rect 1572 79772 1588 79806
rect 122 79686 138 79720
rect 1572 79686 1588 79720
rect 122 79600 138 79634
rect 1572 79600 1588 79634
rect 122 79514 138 79548
rect 1572 79514 1588 79548
rect 122 79428 138 79462
rect 1572 79428 1588 79462
rect 122 79342 138 79376
rect 1572 79342 1588 79376
rect 122 79256 138 79290
rect 1572 79256 1588 79290
rect 122 79170 138 79204
rect 1572 79170 1588 79204
rect 122 79084 138 79118
rect 1572 79084 1588 79118
rect 122 78998 138 79032
rect 1572 78998 1588 79032
rect 122 78912 138 78946
rect 1572 78912 1588 78946
rect 122 78826 138 78860
rect 1572 78826 1588 78860
rect 122 78740 138 78774
rect 1572 78740 1588 78774
rect 122 78654 138 78688
rect 1572 78654 1588 78688
rect 122 78568 138 78602
rect 1572 78568 1588 78602
rect 122 78482 138 78516
rect 1572 78482 1588 78516
rect 122 78396 138 78430
rect 1572 78396 1588 78430
rect 122 78310 138 78344
rect 1572 78310 1588 78344
rect 122 78224 138 78258
rect 1572 78224 1588 78258
rect 122 78138 138 78172
rect 1572 78138 1588 78172
rect 122 78052 138 78086
rect 1572 78052 1588 78086
rect 122 77966 138 78000
rect 1572 77966 1588 78000
rect 122 77880 138 77914
rect 1572 77880 1588 77914
rect 122 77794 138 77828
rect 1572 77794 1588 77828
rect 122 77708 138 77742
rect 1572 77708 1588 77742
rect 122 77622 138 77656
rect 1572 77622 1588 77656
rect 122 77536 138 77570
rect 1572 77536 1588 77570
rect 122 77450 138 77484
rect 1572 77450 1588 77484
rect 122 77364 138 77398
rect 1572 77364 1588 77398
rect 122 77278 138 77312
rect 1572 77278 1588 77312
rect 122 77192 138 77226
rect 1572 77192 1588 77226
rect 122 77106 138 77140
rect 1572 77106 1588 77140
rect 122 77020 138 77054
rect 1572 77020 1588 77054
rect 122 76934 138 76968
rect 1572 76934 1588 76968
rect 122 76848 138 76882
rect 1572 76848 1588 76882
rect 122 76762 138 76796
rect 1572 76762 1588 76796
rect 122 76676 138 76710
rect 1572 76676 1588 76710
rect 122 76590 138 76624
rect 1572 76590 1588 76624
rect 122 76504 138 76538
rect 1572 76504 1588 76538
rect 122 76418 138 76452
rect 1572 76418 1588 76452
rect 122 76332 138 76366
rect 1572 76332 1588 76366
rect 122 76246 138 76280
rect 1572 76246 1588 76280
rect 122 76160 138 76194
rect 1572 76160 1588 76194
rect 122 76074 138 76108
rect 1572 76074 1588 76108
rect 122 75988 138 76022
rect 1572 75988 1588 76022
rect 122 75902 138 75936
rect 1572 75902 1588 75936
rect 122 75816 138 75850
rect 1572 75816 1588 75850
rect 122 75730 138 75764
rect 1572 75730 1588 75764
rect 122 75644 138 75678
rect 1572 75644 1588 75678
rect 122 75558 138 75592
rect 1572 75558 1588 75592
rect 122 75472 138 75506
rect 1572 75472 1588 75506
rect 122 75386 138 75420
rect 1572 75386 1588 75420
rect 122 75300 138 75334
rect 1572 75300 1588 75334
rect 122 75214 138 75248
rect 1572 75214 1588 75248
rect 122 75128 138 75162
rect 1572 75128 1588 75162
rect 122 75042 138 75076
rect 1572 75042 1588 75076
rect 122 74956 138 74990
rect 1572 74956 1588 74990
rect 122 74870 138 74904
rect 1572 74870 1588 74904
rect 122 74784 138 74818
rect 1572 74784 1588 74818
rect 122 74698 138 74732
rect 1572 74698 1588 74732
rect 122 74612 138 74646
rect 1572 74612 1588 74646
rect 122 74526 138 74560
rect 1572 74526 1588 74560
rect 122 74440 138 74474
rect 1572 74440 1588 74474
rect 122 74354 138 74388
rect 1572 74354 1588 74388
rect 122 74268 138 74302
rect 1572 74268 1588 74302
rect 122 74182 138 74216
rect 1572 74182 1588 74216
rect 122 74096 138 74130
rect 1572 74096 1588 74130
rect 122 74010 138 74044
rect 1572 74010 1588 74044
rect 122 73924 138 73958
rect 1572 73924 1588 73958
rect 122 73838 138 73872
rect 1572 73838 1588 73872
rect 122 73752 138 73786
rect 1572 73752 1588 73786
rect 122 73666 138 73700
rect 1572 73666 1588 73700
rect 122 73580 138 73614
rect 1572 73580 1588 73614
rect 122 73494 138 73528
rect 1572 73494 1588 73528
rect 122 73408 138 73442
rect 1572 73408 1588 73442
rect 122 73322 138 73356
rect 1572 73322 1588 73356
rect 122 73236 138 73270
rect 1572 73236 1588 73270
rect 122 73150 138 73184
rect 1572 73150 1588 73184
rect 122 73064 138 73098
rect 1572 73064 1588 73098
rect 122 72978 138 73012
rect 1572 72978 1588 73012
rect 122 72892 138 72926
rect 1572 72892 1588 72926
rect 122 72806 138 72840
rect 1572 72806 1588 72840
rect 122 72720 138 72754
rect 1572 72720 1588 72754
rect 122 72634 138 72668
rect 1572 72634 1588 72668
rect 122 72548 138 72582
rect 1572 72548 1588 72582
rect 122 72462 138 72496
rect 1572 72462 1588 72496
rect 122 72376 138 72410
rect 1572 72376 1588 72410
rect 122 72290 138 72324
rect 1572 72290 1588 72324
rect 122 72204 138 72238
rect 1572 72204 1588 72238
rect 122 72118 138 72152
rect 1572 72118 1588 72152
rect 122 72032 138 72066
rect 1572 72032 1588 72066
rect 122 71946 138 71980
rect 1572 71946 1588 71980
rect 122 71860 138 71894
rect 1572 71860 1588 71894
rect 122 71774 138 71808
rect 1572 71774 1588 71808
rect 122 71688 138 71722
rect 1572 71688 1588 71722
rect 122 71602 138 71636
rect 1572 71602 1588 71636
rect 122 71516 138 71550
rect 1572 71516 1588 71550
rect 122 71430 138 71464
rect 1572 71430 1588 71464
rect 122 71344 138 71378
rect 1572 71344 1588 71378
rect 122 71258 138 71292
rect 1572 71258 1588 71292
rect 122 71172 138 71206
rect 1572 71172 1588 71206
rect 122 71086 138 71120
rect 1572 71086 1588 71120
rect 122 71000 138 71034
rect 1572 71000 1588 71034
rect 122 70914 138 70948
rect 1572 70914 1588 70948
rect 122 70828 138 70862
rect 1572 70828 1588 70862
rect 122 70742 138 70776
rect 1572 70742 1588 70776
rect 122 70656 138 70690
rect 1572 70656 1588 70690
rect 122 70570 138 70604
rect 1572 70570 1588 70604
rect 122 70484 138 70518
rect 1572 70484 1588 70518
rect 122 70398 138 70432
rect 1572 70398 1588 70432
rect 122 70312 138 70346
rect 1572 70312 1588 70346
rect 122 70226 138 70260
rect 1572 70226 1588 70260
rect 122 70140 138 70174
rect 1572 70140 1588 70174
rect 122 70054 138 70088
rect 1572 70054 1588 70088
rect 122 69968 138 70002
rect 1572 69968 1588 70002
rect 122 69882 138 69916
rect 1572 69882 1588 69916
rect 122 69796 138 69830
rect 1572 69796 1588 69830
rect 122 69710 138 69744
rect 1572 69710 1588 69744
rect 122 69624 138 69658
rect 1572 69624 1588 69658
rect 122 69538 138 69572
rect 1572 69538 1588 69572
rect 122 69452 138 69486
rect 1572 69452 1588 69486
rect 122 69366 138 69400
rect 1572 69366 1588 69400
rect 122 69280 138 69314
rect 1572 69280 1588 69314
rect 122 69194 138 69228
rect 1572 69194 1588 69228
rect 122 69108 138 69142
rect 1572 69108 1588 69142
rect 122 69022 138 69056
rect 1572 69022 1588 69056
rect 122 68936 138 68970
rect 1572 68936 1588 68970
rect 122 68850 138 68884
rect 1572 68850 1588 68884
rect 122 68764 138 68798
rect 1572 68764 1588 68798
rect 122 68678 138 68712
rect 1572 68678 1588 68712
rect 122 68592 138 68626
rect 1572 68592 1588 68626
rect 122 68506 138 68540
rect 1572 68506 1588 68540
rect 122 68420 138 68454
rect 1572 68420 1588 68454
rect 122 68334 138 68368
rect 1572 68334 1588 68368
rect 122 68248 138 68282
rect 1572 68248 1588 68282
rect 122 68162 138 68196
rect 1572 68162 1588 68196
rect 122 68076 138 68110
rect 1572 68076 1588 68110
rect 122 67990 138 68024
rect 1572 67990 1588 68024
rect 122 67904 138 67938
rect 1572 67904 1588 67938
rect 122 67818 138 67852
rect 1572 67818 1588 67852
rect 122 67732 138 67766
rect 1572 67732 1588 67766
rect 122 67646 138 67680
rect 1572 67646 1588 67680
rect 122 67560 138 67594
rect 1572 67560 1588 67594
rect 122 67474 138 67508
rect 1572 67474 1588 67508
rect 122 67388 138 67422
rect 1572 67388 1588 67422
rect 122 67302 138 67336
rect 1572 67302 1588 67336
rect 122 67216 138 67250
rect 1572 67216 1588 67250
rect 122 67130 138 67164
rect 1572 67130 1588 67164
rect 122 67044 138 67078
rect 1572 67044 1588 67078
rect 122 66958 138 66992
rect 1572 66958 1588 66992
rect 122 66872 138 66906
rect 1572 66872 1588 66906
rect 122 66786 138 66820
rect 1572 66786 1588 66820
rect 122 66700 138 66734
rect 1572 66700 1588 66734
rect 122 66614 138 66648
rect 1572 66614 1588 66648
rect 122 66528 138 66562
rect 1572 66528 1588 66562
rect 122 66442 138 66476
rect 1572 66442 1588 66476
rect 122 66356 138 66390
rect 1572 66356 1588 66390
rect 122 66270 138 66304
rect 1572 66270 1588 66304
rect 122 66184 138 66218
rect 1572 66184 1588 66218
rect 122 66098 138 66132
rect 1572 66098 1588 66132
rect 122 66012 138 66046
rect 1572 66012 1588 66046
rect 122 65926 138 65960
rect 1572 65926 1588 65960
rect 122 65840 138 65874
rect 1572 65840 1588 65874
rect 122 65754 138 65788
rect 1572 65754 1588 65788
rect 122 65668 138 65702
rect 1572 65668 1588 65702
rect 122 65582 138 65616
rect 1572 65582 1588 65616
rect 122 65496 138 65530
rect 1572 65496 1588 65530
rect 122 65410 138 65444
rect 1572 65410 1588 65444
rect 122 65324 138 65358
rect 1572 65324 1588 65358
rect 122 65238 138 65272
rect 1572 65238 1588 65272
rect 122 65152 138 65186
rect 1572 65152 1588 65186
rect 122 65066 138 65100
rect 1572 65066 1588 65100
rect 122 64980 138 65014
rect 1572 64980 1588 65014
rect 122 64894 138 64928
rect 1572 64894 1588 64928
rect 122 64808 138 64842
rect 1572 64808 1588 64842
rect 122 64722 138 64756
rect 1572 64722 1588 64756
rect 122 64636 138 64670
rect 1572 64636 1588 64670
rect 122 64550 138 64584
rect 1572 64550 1588 64584
rect 122 64464 138 64498
rect 1572 64464 1588 64498
rect 122 64378 138 64412
rect 1572 64378 1588 64412
rect 122 64292 138 64326
rect 1572 64292 1588 64326
rect 122 64206 138 64240
rect 1572 64206 1588 64240
rect 122 64120 138 64154
rect 1572 64120 1588 64154
rect 122 64034 138 64068
rect 1572 64034 1588 64068
rect 122 63948 138 63982
rect 1572 63948 1588 63982
rect 122 63862 138 63896
rect 1572 63862 1588 63896
rect 122 63776 138 63810
rect 1572 63776 1588 63810
rect 122 63690 138 63724
rect 1572 63690 1588 63724
rect 122 63604 138 63638
rect 1572 63604 1588 63638
rect 122 63518 138 63552
rect 1572 63518 1588 63552
rect 122 63432 138 63466
rect 1572 63432 1588 63466
rect 122 63346 138 63380
rect 1572 63346 1588 63380
rect 122 63260 138 63294
rect 1572 63260 1588 63294
rect 122 63174 138 63208
rect 1572 63174 1588 63208
rect 122 63088 138 63122
rect 1572 63088 1588 63122
rect 122 63002 138 63036
rect 1572 63002 1588 63036
rect 122 62916 138 62950
rect 1572 62916 1588 62950
rect 122 62830 138 62864
rect 1572 62830 1588 62864
rect 122 62744 138 62778
rect 1572 62744 1588 62778
rect 122 62658 138 62692
rect 1572 62658 1588 62692
rect 122 62572 138 62606
rect 1572 62572 1588 62606
rect 122 62486 138 62520
rect 1572 62486 1588 62520
rect 122 62400 138 62434
rect 1572 62400 1588 62434
rect 122 62314 138 62348
rect 1572 62314 1588 62348
rect 122 62228 138 62262
rect 1572 62228 1588 62262
rect 122 62142 138 62176
rect 1572 62142 1588 62176
rect 122 62056 138 62090
rect 1572 62056 1588 62090
rect 122 61970 138 62004
rect 1572 61970 1588 62004
rect 122 61884 138 61918
rect 1572 61884 1588 61918
rect 122 61798 138 61832
rect 1572 61798 1588 61832
rect 122 61712 138 61746
rect 1572 61712 1588 61746
rect 122 61626 138 61660
rect 1572 61626 1588 61660
rect 122 61540 138 61574
rect 1572 61540 1588 61574
rect 122 61454 138 61488
rect 1572 61454 1588 61488
rect 122 61368 138 61402
rect 1572 61368 1588 61402
rect 122 61282 138 61316
rect 1572 61282 1588 61316
rect 122 61196 138 61230
rect 1572 61196 1588 61230
rect 122 61110 138 61144
rect 1572 61110 1588 61144
rect 122 61024 138 61058
rect 1572 61024 1588 61058
rect 122 60938 138 60972
rect 1572 60938 1588 60972
rect 122 60852 138 60886
rect 1572 60852 1588 60886
rect 122 60766 138 60800
rect 1572 60766 1588 60800
rect 122 60680 138 60714
rect 1572 60680 1588 60714
rect 122 60594 138 60628
rect 1572 60594 1588 60628
rect 122 60508 138 60542
rect 1572 60508 1588 60542
rect 122 60422 138 60456
rect 1572 60422 1588 60456
rect 122 60336 138 60370
rect 1572 60336 1588 60370
rect 122 60250 138 60284
rect 1572 60250 1588 60284
rect 122 60164 138 60198
rect 1572 60164 1588 60198
rect 122 60078 138 60112
rect 1572 60078 1588 60112
rect 122 59992 138 60026
rect 1572 59992 1588 60026
rect 122 59906 138 59940
rect 1572 59906 1588 59940
rect 122 59820 138 59854
rect 1572 59820 1588 59854
rect 122 59734 138 59768
rect 1572 59734 1588 59768
rect 122 59648 138 59682
rect 1572 59648 1588 59682
rect 122 59562 138 59596
rect 1572 59562 1588 59596
rect 122 59476 138 59510
rect 1572 59476 1588 59510
rect 122 59390 138 59424
rect 1572 59390 1588 59424
rect 122 59304 138 59338
rect 1572 59304 1588 59338
rect 122 59218 138 59252
rect 1572 59218 1588 59252
rect 122 59132 138 59166
rect 1572 59132 1588 59166
rect 122 59046 138 59080
rect 1572 59046 1588 59080
rect 122 58960 138 58994
rect 1572 58960 1588 58994
rect 122 58874 138 58908
rect 1572 58874 1588 58908
rect 122 58788 138 58822
rect 1572 58788 1588 58822
rect 122 58702 138 58736
rect 1572 58702 1588 58736
rect 122 58616 138 58650
rect 1572 58616 1588 58650
rect 122 58530 138 58564
rect 1572 58530 1588 58564
rect 122 58444 138 58478
rect 1572 58444 1588 58478
rect 122 58358 138 58392
rect 1572 58358 1588 58392
rect 122 58272 138 58306
rect 1572 58272 1588 58306
rect 122 58186 138 58220
rect 1572 58186 1588 58220
rect 122 58100 138 58134
rect 1572 58100 1588 58134
rect 122 58014 138 58048
rect 1572 58014 1588 58048
rect 122 57928 138 57962
rect 1572 57928 1588 57962
rect 122 57842 138 57876
rect 1572 57842 1588 57876
rect 122 57756 138 57790
rect 1572 57756 1588 57790
rect 122 57670 138 57704
rect 1572 57670 1588 57704
rect 122 57584 138 57618
rect 1572 57584 1588 57618
rect 122 57498 138 57532
rect 1572 57498 1588 57532
rect 122 57412 138 57446
rect 1572 57412 1588 57446
rect 122 57326 138 57360
rect 1572 57326 1588 57360
rect 122 57240 138 57274
rect 1572 57240 1588 57274
rect 122 57154 138 57188
rect 1572 57154 1588 57188
rect 122 57068 138 57102
rect 1572 57068 1588 57102
rect 122 56982 138 57016
rect 1572 56982 1588 57016
rect 122 56896 138 56930
rect 1572 56896 1588 56930
rect 122 56810 138 56844
rect 1572 56810 1588 56844
rect 122 56724 138 56758
rect 1572 56724 1588 56758
rect 122 56638 138 56672
rect 1572 56638 1588 56672
rect 122 56552 138 56586
rect 1572 56552 1588 56586
rect 122 56466 138 56500
rect 1572 56466 1588 56500
rect 122 56380 138 56414
rect 1572 56380 1588 56414
rect 122 56294 138 56328
rect 1572 56294 1588 56328
rect 122 56208 138 56242
rect 1572 56208 1588 56242
rect 122 56122 138 56156
rect 1572 56122 1588 56156
rect 122 56036 138 56070
rect 1572 56036 1588 56070
rect 122 55950 138 55984
rect 1572 55950 1588 55984
rect 122 55864 138 55898
rect 1572 55864 1588 55898
rect 122 55778 138 55812
rect 1572 55778 1588 55812
rect 122 55692 138 55726
rect 1572 55692 1588 55726
rect 122 55606 138 55640
rect 1572 55606 1588 55640
rect 122 55520 138 55554
rect 1572 55520 1588 55554
rect 122 55434 138 55468
rect 1572 55434 1588 55468
rect 122 55348 138 55382
rect 1572 55348 1588 55382
rect 122 55262 138 55296
rect 1572 55262 1588 55296
rect 122 55176 138 55210
rect 1572 55176 1588 55210
rect 122 55090 138 55124
rect 1572 55090 1588 55124
rect 122 55004 138 55038
rect 1572 55004 1588 55038
rect 122 54918 138 54952
rect 1572 54918 1588 54952
rect 122 54832 138 54866
rect 1572 54832 1588 54866
rect 122 54746 138 54780
rect 1572 54746 1588 54780
rect 122 54660 138 54694
rect 1572 54660 1588 54694
rect 122 54574 138 54608
rect 1572 54574 1588 54608
rect 122 54488 138 54522
rect 1572 54488 1588 54522
rect 122 54402 138 54436
rect 1572 54402 1588 54436
rect 122 54316 138 54350
rect 1572 54316 1588 54350
rect 122 54230 138 54264
rect 1572 54230 1588 54264
rect 122 54144 138 54178
rect 1572 54144 1588 54178
rect 122 54058 138 54092
rect 1572 54058 1588 54092
rect 122 53972 138 54006
rect 1572 53972 1588 54006
rect 122 53886 138 53920
rect 1572 53886 1588 53920
rect 122 53800 138 53834
rect 1572 53800 1588 53834
rect 122 53714 138 53748
rect 1572 53714 1588 53748
rect 122 53628 138 53662
rect 1572 53628 1588 53662
rect 122 53542 138 53576
rect 1572 53542 1588 53576
rect 122 53456 138 53490
rect 1572 53456 1588 53490
rect 122 53370 138 53404
rect 1572 53370 1588 53404
rect 122 53284 138 53318
rect 1572 53284 1588 53318
rect 122 53198 138 53232
rect 1572 53198 1588 53232
rect 122 53112 138 53146
rect 1572 53112 1588 53146
rect 122 53026 138 53060
rect 1572 53026 1588 53060
rect 122 52940 138 52974
rect 1572 52940 1588 52974
rect 122 52854 138 52888
rect 1572 52854 1588 52888
rect 122 52768 138 52802
rect 1572 52768 1588 52802
rect 122 52682 138 52716
rect 1572 52682 1588 52716
rect 122 52596 138 52630
rect 1572 52596 1588 52630
rect 122 52510 138 52544
rect 1572 52510 1588 52544
rect 122 52424 138 52458
rect 1572 52424 1588 52458
rect 122 52338 138 52372
rect 1572 52338 1588 52372
rect 122 52252 138 52286
rect 1572 52252 1588 52286
rect 122 52166 138 52200
rect 1572 52166 1588 52200
rect 122 52080 138 52114
rect 1572 52080 1588 52114
rect 122 51994 138 52028
rect 1572 51994 1588 52028
rect 122 51908 138 51942
rect 1572 51908 1588 51942
rect 122 51822 138 51856
rect 1572 51822 1588 51856
rect 122 51736 138 51770
rect 1572 51736 1588 51770
rect 122 51650 138 51684
rect 1572 51650 1588 51684
rect 122 51564 138 51598
rect 1572 51564 1588 51598
rect 122 51478 138 51512
rect 1572 51478 1588 51512
rect 122 51392 138 51426
rect 1572 51392 1588 51426
rect 122 51306 138 51340
rect 1572 51306 1588 51340
rect 122 51220 138 51254
rect 1572 51220 1588 51254
rect 122 51134 138 51168
rect 1572 51134 1588 51168
rect 122 51048 138 51082
rect 1572 51048 1588 51082
rect 122 50962 138 50996
rect 1572 50962 1588 50996
rect 122 50876 138 50910
rect 1572 50876 1588 50910
rect 122 50790 138 50824
rect 1572 50790 1588 50824
rect 122 50704 138 50738
rect 1572 50704 1588 50738
rect 122 50618 138 50652
rect 1572 50618 1588 50652
rect 122 50532 138 50566
rect 1572 50532 1588 50566
rect 122 50446 138 50480
rect 1572 50446 1588 50480
rect 122 50360 138 50394
rect 1572 50360 1588 50394
rect 122 50274 138 50308
rect 1572 50274 1588 50308
rect 122 50188 138 50222
rect 1572 50188 1588 50222
rect 122 50102 138 50136
rect 1572 50102 1588 50136
rect 122 50016 138 50050
rect 1572 50016 1588 50050
rect 122 49930 138 49964
rect 1572 49930 1588 49964
rect 122 49844 138 49878
rect 1572 49844 1588 49878
rect 122 49758 138 49792
rect 1572 49758 1588 49792
rect 122 49672 138 49706
rect 1572 49672 1588 49706
rect 122 49586 138 49620
rect 1572 49586 1588 49620
rect 122 49500 138 49534
rect 1572 49500 1588 49534
rect 122 49414 138 49448
rect 1572 49414 1588 49448
rect 122 49328 138 49362
rect 1572 49328 1588 49362
rect 122 49242 138 49276
rect 1572 49242 1588 49276
rect 122 49156 138 49190
rect 1572 49156 1588 49190
rect 122 49070 138 49104
rect 1572 49070 1588 49104
rect 122 48984 138 49018
rect 1572 48984 1588 49018
rect 122 48898 138 48932
rect 1572 48898 1588 48932
rect 122 48812 138 48846
rect 1572 48812 1588 48846
rect 122 48726 138 48760
rect 1572 48726 1588 48760
rect 122 48640 138 48674
rect 1572 48640 1588 48674
rect 122 48554 138 48588
rect 1572 48554 1588 48588
rect 122 48468 138 48502
rect 1572 48468 1588 48502
rect 122 48382 138 48416
rect 1572 48382 1588 48416
rect 122 48296 138 48330
rect 1572 48296 1588 48330
rect 122 48210 138 48244
rect 1572 48210 1588 48244
rect 122 48124 138 48158
rect 1572 48124 1588 48158
rect 122 48038 138 48072
rect 1572 48038 1588 48072
rect 122 47952 138 47986
rect 1572 47952 1588 47986
rect 122 47866 138 47900
rect 1572 47866 1588 47900
rect 122 47780 138 47814
rect 1572 47780 1588 47814
rect 122 47694 138 47728
rect 1572 47694 1588 47728
rect 122 47608 138 47642
rect 1572 47608 1588 47642
rect 122 47522 138 47556
rect 1572 47522 1588 47556
rect 122 47436 138 47470
rect 1572 47436 1588 47470
rect 122 47350 138 47384
rect 1572 47350 1588 47384
rect 122 47264 138 47298
rect 1572 47264 1588 47298
rect 122 47178 138 47212
rect 1572 47178 1588 47212
rect 122 47092 138 47126
rect 1572 47092 1588 47126
rect 122 47006 138 47040
rect 1572 47006 1588 47040
rect 122 46920 138 46954
rect 1572 46920 1588 46954
rect 122 46834 138 46868
rect 1572 46834 1588 46868
rect 122 46748 138 46782
rect 1572 46748 1588 46782
rect 122 46662 138 46696
rect 1572 46662 1588 46696
rect 122 46576 138 46610
rect 1572 46576 1588 46610
rect 122 46490 138 46524
rect 1572 46490 1588 46524
rect 122 46404 138 46438
rect 1572 46404 1588 46438
rect 122 46318 138 46352
rect 1572 46318 1588 46352
rect 122 46232 138 46266
rect 1572 46232 1588 46266
rect 122 46146 138 46180
rect 1572 46146 1588 46180
rect 122 46060 138 46094
rect 1572 46060 1588 46094
rect 122 45974 138 46008
rect 1572 45974 1588 46008
rect 122 45888 138 45922
rect 1572 45888 1588 45922
rect 122 45802 138 45836
rect 1572 45802 1588 45836
rect 122 45716 138 45750
rect 1572 45716 1588 45750
rect 122 45630 138 45664
rect 1572 45630 1588 45664
rect 122 45544 138 45578
rect 1572 45544 1588 45578
rect 122 45458 138 45492
rect 1572 45458 1588 45492
rect 122 45372 138 45406
rect 1572 45372 1588 45406
rect 122 45286 138 45320
rect 1572 45286 1588 45320
rect 122 45200 138 45234
rect 1572 45200 1588 45234
rect 122 45114 138 45148
rect 1572 45114 1588 45148
rect 122 45028 138 45062
rect 1572 45028 1588 45062
rect 122 44942 138 44976
rect 1572 44942 1588 44976
rect 122 44856 138 44890
rect 1572 44856 1588 44890
rect 122 44770 138 44804
rect 1572 44770 1588 44804
rect 122 44684 138 44718
rect 1572 44684 1588 44718
rect 122 44598 138 44632
rect 1572 44598 1588 44632
rect 122 44512 138 44546
rect 1572 44512 1588 44546
rect 122 44426 138 44460
rect 1572 44426 1588 44460
rect 122 44340 138 44374
rect 1572 44340 1588 44374
rect 122 44254 138 44288
rect 1572 44254 1588 44288
rect 122 44168 138 44202
rect 1572 44168 1588 44202
rect 122 44082 138 44116
rect 1572 44082 1588 44116
rect 122 43996 138 44030
rect 1572 43996 1588 44030
rect 122 43910 138 43944
rect 1572 43910 1588 43944
rect 122 43824 138 43858
rect 1572 43824 1588 43858
rect 122 43738 138 43772
rect 1572 43738 1588 43772
rect 122 43652 138 43686
rect 1572 43652 1588 43686
rect 122 43566 138 43600
rect 1572 43566 1588 43600
rect 122 43480 138 43514
rect 1572 43480 1588 43514
rect 122 43394 138 43428
rect 1572 43394 1588 43428
rect 122 43308 138 43342
rect 1572 43308 1588 43342
rect 122 43222 138 43256
rect 1572 43222 1588 43256
rect 122 43136 138 43170
rect 1572 43136 1588 43170
rect 122 43050 138 43084
rect 1572 43050 1588 43084
rect 122 42964 138 42998
rect 1572 42964 1588 42998
rect 122 42878 138 42912
rect 1572 42878 1588 42912
rect 122 42792 138 42826
rect 1572 42792 1588 42826
rect 122 42706 138 42740
rect 1572 42706 1588 42740
rect 122 42620 138 42654
rect 1572 42620 1588 42654
rect 122 42534 138 42568
rect 1572 42534 1588 42568
rect 122 42448 138 42482
rect 1572 42448 1588 42482
rect 122 42362 138 42396
rect 1572 42362 1588 42396
rect 122 42276 138 42310
rect 1572 42276 1588 42310
rect 122 42190 138 42224
rect 1572 42190 1588 42224
rect 122 42104 138 42138
rect 1572 42104 1588 42138
rect 122 42018 138 42052
rect 1572 42018 1588 42052
rect 122 41932 138 41966
rect 1572 41932 1588 41966
rect 122 41846 138 41880
rect 1572 41846 1588 41880
rect 122 41760 138 41794
rect 1572 41760 1588 41794
rect 122 41674 138 41708
rect 1572 41674 1588 41708
rect 122 41588 138 41622
rect 1572 41588 1588 41622
rect 122 41502 138 41536
rect 1572 41502 1588 41536
rect 122 41416 138 41450
rect 1572 41416 1588 41450
rect 122 41330 138 41364
rect 1572 41330 1588 41364
rect 122 41244 138 41278
rect 1572 41244 1588 41278
rect 122 41158 138 41192
rect 1572 41158 1588 41192
rect 122 41072 138 41106
rect 1572 41072 1588 41106
rect 122 40986 138 41020
rect 1572 40986 1588 41020
rect 122 40900 138 40934
rect 1572 40900 1588 40934
rect 122 40814 138 40848
rect 1572 40814 1588 40848
rect 122 40728 138 40762
rect 1572 40728 1588 40762
rect 122 40642 138 40676
rect 1572 40642 1588 40676
rect 122 40556 138 40590
rect 1572 40556 1588 40590
rect 122 40470 138 40504
rect 1572 40470 1588 40504
rect 122 40384 138 40418
rect 1572 40384 1588 40418
rect 122 40298 138 40332
rect 1572 40298 1588 40332
rect 122 40212 138 40246
rect 1572 40212 1588 40246
rect 122 40126 138 40160
rect 1572 40126 1588 40160
rect 122 40040 138 40074
rect 1572 40040 1588 40074
rect 122 39954 138 39988
rect 1572 39954 1588 39988
rect 122 39868 138 39902
rect 1572 39868 1588 39902
rect 122 39782 138 39816
rect 1572 39782 1588 39816
rect 122 39696 138 39730
rect 1572 39696 1588 39730
rect 122 39610 138 39644
rect 1572 39610 1588 39644
rect 122 39524 138 39558
rect 1572 39524 1588 39558
rect 122 39438 138 39472
rect 1572 39438 1588 39472
rect 122 39352 138 39386
rect 1572 39352 1588 39386
rect 122 39266 138 39300
rect 1572 39266 1588 39300
rect 122 39180 138 39214
rect 1572 39180 1588 39214
rect 122 39094 138 39128
rect 1572 39094 1588 39128
rect 122 39008 138 39042
rect 1572 39008 1588 39042
rect 122 38922 138 38956
rect 1572 38922 1588 38956
rect 122 38836 138 38870
rect 1572 38836 1588 38870
rect 122 38750 138 38784
rect 1572 38750 1588 38784
rect 122 38664 138 38698
rect 1572 38664 1588 38698
rect 122 38578 138 38612
rect 1572 38578 1588 38612
rect 122 38492 138 38526
rect 1572 38492 1588 38526
rect 122 38406 138 38440
rect 1572 38406 1588 38440
rect 122 38320 138 38354
rect 1572 38320 1588 38354
rect 122 38234 138 38268
rect 1572 38234 1588 38268
rect 122 38148 138 38182
rect 1572 38148 1588 38182
rect 122 38062 138 38096
rect 1572 38062 1588 38096
rect 122 37976 138 38010
rect 1572 37976 1588 38010
rect 122 37890 138 37924
rect 1572 37890 1588 37924
rect 122 37804 138 37838
rect 1572 37804 1588 37838
rect 122 37718 138 37752
rect 1572 37718 1588 37752
rect 122 37632 138 37666
rect 1572 37632 1588 37666
rect 122 37546 138 37580
rect 1572 37546 1588 37580
rect 122 37460 138 37494
rect 1572 37460 1588 37494
rect 122 37374 138 37408
rect 1572 37374 1588 37408
rect 122 37288 138 37322
rect 1572 37288 1588 37322
rect 122 37202 138 37236
rect 1572 37202 1588 37236
rect 122 37116 138 37150
rect 1572 37116 1588 37150
rect 122 37030 138 37064
rect 1572 37030 1588 37064
rect 122 36944 138 36978
rect 1572 36944 1588 36978
rect 122 36858 138 36892
rect 1572 36858 1588 36892
rect 122 36772 138 36806
rect 1572 36772 1588 36806
rect 122 36686 138 36720
rect 1572 36686 1588 36720
rect 122 36600 138 36634
rect 1572 36600 1588 36634
rect 122 36514 138 36548
rect 1572 36514 1588 36548
rect 122 36428 138 36462
rect 1572 36428 1588 36462
rect 122 36342 138 36376
rect 1572 36342 1588 36376
rect 122 36256 138 36290
rect 1572 36256 1588 36290
rect 122 36170 138 36204
rect 1572 36170 1588 36204
rect 122 36084 138 36118
rect 1572 36084 1588 36118
rect 122 35998 138 36032
rect 1572 35998 1588 36032
rect 122 35912 138 35946
rect 1572 35912 1588 35946
rect 122 35826 138 35860
rect 1572 35826 1588 35860
rect 122 35740 138 35774
rect 1572 35740 1588 35774
rect 122 35654 138 35688
rect 1572 35654 1588 35688
rect 122 35568 138 35602
rect 1572 35568 1588 35602
rect 122 35482 138 35516
rect 1572 35482 1588 35516
rect 122 35396 138 35430
rect 1572 35396 1588 35430
rect 122 35310 138 35344
rect 1572 35310 1588 35344
rect 122 35224 138 35258
rect 1572 35224 1588 35258
rect 122 35138 138 35172
rect 1572 35138 1588 35172
rect 122 35052 138 35086
rect 1572 35052 1588 35086
rect 122 34966 138 35000
rect 1572 34966 1588 35000
rect 122 34880 138 34914
rect 1572 34880 1588 34914
rect 122 34794 138 34828
rect 1572 34794 1588 34828
rect 122 34708 138 34742
rect 1572 34708 1588 34742
rect 122 34622 138 34656
rect 1572 34622 1588 34656
rect 122 34536 138 34570
rect 1572 34536 1588 34570
rect 122 34450 138 34484
rect 1572 34450 1588 34484
rect 122 34364 138 34398
rect 1572 34364 1588 34398
rect 122 34278 138 34312
rect 1572 34278 1588 34312
rect 122 34192 138 34226
rect 1572 34192 1588 34226
rect 122 34106 138 34140
rect 1572 34106 1588 34140
rect 122 34020 138 34054
rect 1572 34020 1588 34054
rect 122 33934 138 33968
rect 1572 33934 1588 33968
rect 122 33848 138 33882
rect 1572 33848 1588 33882
rect 122 33762 138 33796
rect 1572 33762 1588 33796
rect 122 33676 138 33710
rect 1572 33676 1588 33710
rect 122 33590 138 33624
rect 1572 33590 1588 33624
rect 122 33504 138 33538
rect 1572 33504 1588 33538
rect 122 33418 138 33452
rect 1572 33418 1588 33452
rect 122 33332 138 33366
rect 1572 33332 1588 33366
rect 122 33246 138 33280
rect 1572 33246 1588 33280
rect 122 33160 138 33194
rect 1572 33160 1588 33194
rect 122 33074 138 33108
rect 1572 33074 1588 33108
rect 122 32988 138 33022
rect 1572 32988 1588 33022
rect 122 32902 138 32936
rect 1572 32902 1588 32936
rect 122 32816 138 32850
rect 1572 32816 1588 32850
rect 122 32730 138 32764
rect 1572 32730 1588 32764
rect 122 32644 138 32678
rect 1572 32644 1588 32678
rect 122 32558 138 32592
rect 1572 32558 1588 32592
rect 122 32472 138 32506
rect 1572 32472 1588 32506
rect 122 32386 138 32420
rect 1572 32386 1588 32420
rect 122 32300 138 32334
rect 1572 32300 1588 32334
rect 122 32214 138 32248
rect 1572 32214 1588 32248
rect 122 32128 138 32162
rect 1572 32128 1588 32162
rect 122 32042 138 32076
rect 1572 32042 1588 32076
rect 122 31956 138 31990
rect 1572 31956 1588 31990
rect 122 31870 138 31904
rect 1572 31870 1588 31904
rect 122 31784 138 31818
rect 1572 31784 1588 31818
rect 122 31698 138 31732
rect 1572 31698 1588 31732
rect 122 31612 138 31646
rect 1572 31612 1588 31646
rect 122 31526 138 31560
rect 1572 31526 1588 31560
rect 122 31440 138 31474
rect 1572 31440 1588 31474
rect 122 31354 138 31388
rect 1572 31354 1588 31388
rect 122 31268 138 31302
rect 1572 31268 1588 31302
rect 122 31182 138 31216
rect 1572 31182 1588 31216
rect 122 31096 138 31130
rect 1572 31096 1588 31130
rect 122 31010 138 31044
rect 1572 31010 1588 31044
rect 122 30924 138 30958
rect 1572 30924 1588 30958
rect 122 30838 138 30872
rect 1572 30838 1588 30872
rect 122 30752 138 30786
rect 1572 30752 1588 30786
rect 122 30666 138 30700
rect 1572 30666 1588 30700
rect 122 30580 138 30614
rect 1572 30580 1588 30614
rect 122 30494 138 30528
rect 1572 30494 1588 30528
rect 122 30408 138 30442
rect 1572 30408 1588 30442
rect 122 30322 138 30356
rect 1572 30322 1588 30356
rect 122 30236 138 30270
rect 1572 30236 1588 30270
rect 122 30150 138 30184
rect 1572 30150 1588 30184
rect 122 30064 138 30098
rect 1572 30064 1588 30098
rect 122 29978 138 30012
rect 1572 29978 1588 30012
rect 122 29892 138 29926
rect 1572 29892 1588 29926
rect 122 29806 138 29840
rect 1572 29806 1588 29840
rect 122 29720 138 29754
rect 1572 29720 1588 29754
rect 122 29634 138 29668
rect 1572 29634 1588 29668
rect 122 29548 138 29582
rect 1572 29548 1588 29582
rect 122 29462 138 29496
rect 1572 29462 1588 29496
rect 122 29376 138 29410
rect 1572 29376 1588 29410
rect 122 29290 138 29324
rect 1572 29290 1588 29324
rect 122 29204 138 29238
rect 1572 29204 1588 29238
rect 122 29118 138 29152
rect 1572 29118 1588 29152
rect 122 29032 138 29066
rect 1572 29032 1588 29066
rect 122 28946 138 28980
rect 1572 28946 1588 28980
rect 122 28860 138 28894
rect 1572 28860 1588 28894
rect 122 28774 138 28808
rect 1572 28774 1588 28808
rect 122 28688 138 28722
rect 1572 28688 1588 28722
rect 122 28602 138 28636
rect 1572 28602 1588 28636
rect 122 28516 138 28550
rect 1572 28516 1588 28550
rect 122 28430 138 28464
rect 1572 28430 1588 28464
rect 122 28344 138 28378
rect 1572 28344 1588 28378
rect 122 28258 138 28292
rect 1572 28258 1588 28292
rect 122 28172 138 28206
rect 1572 28172 1588 28206
rect 122 28086 138 28120
rect 1572 28086 1588 28120
rect 122 28000 138 28034
rect 1572 28000 1588 28034
rect 122 27914 138 27948
rect 1572 27914 1588 27948
rect 122 27828 138 27862
rect 1572 27828 1588 27862
rect 122 27742 138 27776
rect 1572 27742 1588 27776
rect 122 27656 138 27690
rect 1572 27656 1588 27690
rect 122 27570 138 27604
rect 1572 27570 1588 27604
rect 122 27484 138 27518
rect 1572 27484 1588 27518
rect 122 27398 138 27432
rect 1572 27398 1588 27432
rect 122 27312 138 27346
rect 1572 27312 1588 27346
rect 122 27226 138 27260
rect 1572 27226 1588 27260
rect 122 27140 138 27174
rect 1572 27140 1588 27174
rect 122 27054 138 27088
rect 1572 27054 1588 27088
rect 122 26968 138 27002
rect 1572 26968 1588 27002
rect 122 26882 138 26916
rect 1572 26882 1588 26916
rect 122 26796 138 26830
rect 1572 26796 1588 26830
rect 122 26710 138 26744
rect 1572 26710 1588 26744
rect 122 26624 138 26658
rect 1572 26624 1588 26658
rect 122 26538 138 26572
rect 1572 26538 1588 26572
rect 122 26452 138 26486
rect 1572 26452 1588 26486
rect 122 26366 138 26400
rect 1572 26366 1588 26400
rect 122 26280 138 26314
rect 1572 26280 1588 26314
rect 122 26194 138 26228
rect 1572 26194 1588 26228
rect 122 26108 138 26142
rect 1572 26108 1588 26142
rect 122 26022 138 26056
rect 1572 26022 1588 26056
rect 122 25936 138 25970
rect 1572 25936 1588 25970
rect 122 25850 138 25884
rect 1572 25850 1588 25884
rect 122 25764 138 25798
rect 1572 25764 1588 25798
rect 122 25678 138 25712
rect 1572 25678 1588 25712
rect 122 25592 138 25626
rect 1572 25592 1588 25626
rect 122 25506 138 25540
rect 1572 25506 1588 25540
rect 122 25420 138 25454
rect 1572 25420 1588 25454
rect 122 25334 138 25368
rect 1572 25334 1588 25368
rect 122 25248 138 25282
rect 1572 25248 1588 25282
rect 122 25162 138 25196
rect 1572 25162 1588 25196
rect 122 25076 138 25110
rect 1572 25076 1588 25110
rect 122 24990 138 25024
rect 1572 24990 1588 25024
rect 122 24904 138 24938
rect 1572 24904 1588 24938
rect 122 24818 138 24852
rect 1572 24818 1588 24852
rect 122 24732 138 24766
rect 1572 24732 1588 24766
rect 122 24646 138 24680
rect 1572 24646 1588 24680
rect 122 24560 138 24594
rect 1572 24560 1588 24594
rect 122 24474 138 24508
rect 1572 24474 1588 24508
rect 122 24388 138 24422
rect 1572 24388 1588 24422
rect 122 24302 138 24336
rect 1572 24302 1588 24336
rect 122 24216 138 24250
rect 1572 24216 1588 24250
rect 122 24130 138 24164
rect 1572 24130 1588 24164
rect 122 24044 138 24078
rect 1572 24044 1588 24078
rect 122 23958 138 23992
rect 1572 23958 1588 23992
rect 122 23872 138 23906
rect 1572 23872 1588 23906
rect 122 23786 138 23820
rect 1572 23786 1588 23820
rect 122 23700 138 23734
rect 1572 23700 1588 23734
rect 122 23614 138 23648
rect 1572 23614 1588 23648
rect 122 23528 138 23562
rect 1572 23528 1588 23562
rect 122 23442 138 23476
rect 1572 23442 1588 23476
rect 122 23356 138 23390
rect 1572 23356 1588 23390
rect 122 23270 138 23304
rect 1572 23270 1588 23304
rect 122 23184 138 23218
rect 1572 23184 1588 23218
rect 122 23098 138 23132
rect 1572 23098 1588 23132
rect 122 23012 138 23046
rect 1572 23012 1588 23046
rect 122 22926 138 22960
rect 1572 22926 1588 22960
rect 122 22840 138 22874
rect 1572 22840 1588 22874
rect 122 22754 138 22788
rect 1572 22754 1588 22788
rect 122 22668 138 22702
rect 1572 22668 1588 22702
rect 122 22582 138 22616
rect 1572 22582 1588 22616
rect 122 22496 138 22530
rect 1572 22496 1588 22530
rect 122 22410 138 22444
rect 1572 22410 1588 22444
rect 122 22324 138 22358
rect 1572 22324 1588 22358
rect 122 22238 138 22272
rect 1572 22238 1588 22272
rect 122 22152 138 22186
rect 1572 22152 1588 22186
rect 122 22066 138 22100
rect 1572 22066 1588 22100
rect 122 21980 138 22014
rect 1572 21980 1588 22014
rect 122 21894 138 21928
rect 1572 21894 1588 21928
rect 122 21808 138 21842
rect 1572 21808 1588 21842
rect 122 21722 138 21756
rect 1572 21722 1588 21756
rect 122 21636 138 21670
rect 1572 21636 1588 21670
rect 122 21550 138 21584
rect 1572 21550 1588 21584
rect 122 21464 138 21498
rect 1572 21464 1588 21498
rect 122 21378 138 21412
rect 1572 21378 1588 21412
rect 122 21292 138 21326
rect 1572 21292 1588 21326
rect 122 21206 138 21240
rect 1572 21206 1588 21240
rect 122 21120 138 21154
rect 1572 21120 1588 21154
rect 122 21034 138 21068
rect 1572 21034 1588 21068
rect 122 20948 138 20982
rect 1572 20948 1588 20982
rect 122 20862 138 20896
rect 1572 20862 1588 20896
rect 122 20776 138 20810
rect 1572 20776 1588 20810
rect 122 20690 138 20724
rect 1572 20690 1588 20724
rect 122 20604 138 20638
rect 1572 20604 1588 20638
rect 122 20518 138 20552
rect 1572 20518 1588 20552
rect 122 20432 138 20466
rect 1572 20432 1588 20466
rect 122 20346 138 20380
rect 1572 20346 1588 20380
rect 122 20260 138 20294
rect 1572 20260 1588 20294
rect 122 20174 138 20208
rect 1572 20174 1588 20208
rect 122 20088 138 20122
rect 1572 20088 1588 20122
rect 122 20002 138 20036
rect 1572 20002 1588 20036
rect 122 19916 138 19950
rect 1572 19916 1588 19950
rect 122 19830 138 19864
rect 1572 19830 1588 19864
rect 122 19744 138 19778
rect 1572 19744 1588 19778
rect 122 19658 138 19692
rect 1572 19658 1588 19692
rect 122 19572 138 19606
rect 1572 19572 1588 19606
rect 122 19486 138 19520
rect 1572 19486 1588 19520
rect 122 19400 138 19434
rect 1572 19400 1588 19434
rect 122 19314 138 19348
rect 1572 19314 1588 19348
rect 122 19228 138 19262
rect 1572 19228 1588 19262
rect 122 19142 138 19176
rect 1572 19142 1588 19176
rect 122 19056 138 19090
rect 1572 19056 1588 19090
rect 122 18970 138 19004
rect 1572 18970 1588 19004
rect 122 18884 138 18918
rect 1572 18884 1588 18918
rect 122 18798 138 18832
rect 1572 18798 1588 18832
rect 122 18712 138 18746
rect 1572 18712 1588 18746
rect 122 18626 138 18660
rect 1572 18626 1588 18660
rect 122 18540 138 18574
rect 1572 18540 1588 18574
rect 122 18454 138 18488
rect 1572 18454 1588 18488
rect 122 18368 138 18402
rect 1572 18368 1588 18402
rect 122 18282 138 18316
rect 1572 18282 1588 18316
rect 122 18196 138 18230
rect 1572 18196 1588 18230
rect 122 18110 138 18144
rect 1572 18110 1588 18144
rect 122 18024 138 18058
rect 1572 18024 1588 18058
rect 122 17938 138 17972
rect 1572 17938 1588 17972
rect 122 17852 138 17886
rect 1572 17852 1588 17886
rect 122 17766 138 17800
rect 1572 17766 1588 17800
rect 122 17680 138 17714
rect 1572 17680 1588 17714
rect 122 17594 138 17628
rect 1572 17594 1588 17628
rect 122 17508 138 17542
rect 1572 17508 1588 17542
rect 122 17422 138 17456
rect 1572 17422 1588 17456
rect 122 17336 138 17370
rect 1572 17336 1588 17370
rect 122 17250 138 17284
rect 1572 17250 1588 17284
rect 122 17164 138 17198
rect 1572 17164 1588 17198
rect 122 17078 138 17112
rect 1572 17078 1588 17112
rect 122 16992 138 17026
rect 1572 16992 1588 17026
rect 122 16906 138 16940
rect 1572 16906 1588 16940
rect 122 16820 138 16854
rect 1572 16820 1588 16854
rect 122 16734 138 16768
rect 1572 16734 1588 16768
rect 122 16648 138 16682
rect 1572 16648 1588 16682
rect 122 16562 138 16596
rect 1572 16562 1588 16596
rect 122 16476 138 16510
rect 1572 16476 1588 16510
rect 122 16390 138 16424
rect 1572 16390 1588 16424
rect 122 16304 138 16338
rect 1572 16304 1588 16338
rect 122 16218 138 16252
rect 1572 16218 1588 16252
rect 122 16132 138 16166
rect 1572 16132 1588 16166
rect 122 16046 138 16080
rect 1572 16046 1588 16080
rect 122 15960 138 15994
rect 1572 15960 1588 15994
rect 122 15874 138 15908
rect 1572 15874 1588 15908
rect 122 15788 138 15822
rect 1572 15788 1588 15822
rect 122 15702 138 15736
rect 1572 15702 1588 15736
rect 122 15616 138 15650
rect 1572 15616 1588 15650
rect 122 15530 138 15564
rect 1572 15530 1588 15564
rect 122 15444 138 15478
rect 1572 15444 1588 15478
rect 122 15358 138 15392
rect 1572 15358 1588 15392
rect 122 15272 138 15306
rect 1572 15272 1588 15306
rect 122 15186 138 15220
rect 1572 15186 1588 15220
rect 122 15100 138 15134
rect 1572 15100 1588 15134
rect 122 15014 138 15048
rect 1572 15014 1588 15048
rect 122 14928 138 14962
rect 1572 14928 1588 14962
rect 122 14842 138 14876
rect 1572 14842 1588 14876
rect 122 14756 138 14790
rect 1572 14756 1588 14790
rect 122 14670 138 14704
rect 1572 14670 1588 14704
rect 122 14584 138 14618
rect 1572 14584 1588 14618
rect 122 14498 138 14532
rect 1572 14498 1588 14532
rect 122 14412 138 14446
rect 1572 14412 1588 14446
rect 122 14326 138 14360
rect 1572 14326 1588 14360
rect 122 14240 138 14274
rect 1572 14240 1588 14274
rect 122 14154 138 14188
rect 1572 14154 1588 14188
rect 122 14068 138 14102
rect 1572 14068 1588 14102
rect 122 13982 138 14016
rect 1572 13982 1588 14016
rect 122 13896 138 13930
rect 1572 13896 1588 13930
rect 122 13810 138 13844
rect 1572 13810 1588 13844
rect 122 13724 138 13758
rect 1572 13724 1588 13758
rect 122 13638 138 13672
rect 1572 13638 1588 13672
rect 122 13552 138 13586
rect 1572 13552 1588 13586
rect 122 13466 138 13500
rect 1572 13466 1588 13500
rect 122 13380 138 13414
rect 1572 13380 1588 13414
rect 122 13294 138 13328
rect 1572 13294 1588 13328
rect 122 13208 138 13242
rect 1572 13208 1588 13242
rect 122 13122 138 13156
rect 1572 13122 1588 13156
rect 122 13036 138 13070
rect 1572 13036 1588 13070
rect 122 12950 138 12984
rect 1572 12950 1588 12984
rect 122 12864 138 12898
rect 1572 12864 1588 12898
rect 122 12778 138 12812
rect 1572 12778 1588 12812
rect 122 12692 138 12726
rect 1572 12692 1588 12726
rect 122 12606 138 12640
rect 1572 12606 1588 12640
rect 122 12520 138 12554
rect 1572 12520 1588 12554
rect 122 12434 138 12468
rect 1572 12434 1588 12468
rect 122 12348 138 12382
rect 1572 12348 1588 12382
rect 122 12262 138 12296
rect 1572 12262 1588 12296
rect 122 12176 138 12210
rect 1572 12176 1588 12210
rect 122 12090 138 12124
rect 1572 12090 1588 12124
rect 122 12004 138 12038
rect 1572 12004 1588 12038
rect 122 11918 138 11952
rect 1572 11918 1588 11952
rect 122 11832 138 11866
rect 1572 11832 1588 11866
rect 122 11746 138 11780
rect 1572 11746 1588 11780
rect 122 11660 138 11694
rect 1572 11660 1588 11694
rect 122 11574 138 11608
rect 1572 11574 1588 11608
rect 122 11488 138 11522
rect 1572 11488 1588 11522
rect 122 11402 138 11436
rect 1572 11402 1588 11436
rect 122 11316 138 11350
rect 1572 11316 1588 11350
rect 122 11230 138 11264
rect 1572 11230 1588 11264
rect 122 11144 138 11178
rect 1572 11144 1588 11178
rect 122 11058 138 11092
rect 1572 11058 1588 11092
rect 122 10972 138 11006
rect 1572 10972 1588 11006
rect 122 10886 138 10920
rect 1572 10886 1588 10920
rect 122 10800 138 10834
rect 1572 10800 1588 10834
rect 122 10714 138 10748
rect 1572 10714 1588 10748
rect 122 10628 138 10662
rect 1572 10628 1588 10662
rect 122 10542 138 10576
rect 1572 10542 1588 10576
rect 122 10456 138 10490
rect 1572 10456 1588 10490
rect 122 10370 138 10404
rect 1572 10370 1588 10404
rect 122 10284 138 10318
rect 1572 10284 1588 10318
rect 122 10198 138 10232
rect 1572 10198 1588 10232
rect 122 10112 138 10146
rect 1572 10112 1588 10146
rect 122 10026 138 10060
rect 1572 10026 1588 10060
rect 122 9940 138 9974
rect 1572 9940 1588 9974
rect 122 9854 138 9888
rect 1572 9854 1588 9888
rect 122 9768 138 9802
rect 1572 9768 1588 9802
rect 122 9682 138 9716
rect 1572 9682 1588 9716
rect 122 9596 138 9630
rect 1572 9596 1588 9630
rect 122 9510 138 9544
rect 1572 9510 1588 9544
rect 122 9424 138 9458
rect 1572 9424 1588 9458
rect 122 9338 138 9372
rect 1572 9338 1588 9372
rect 122 9252 138 9286
rect 1572 9252 1588 9286
rect 122 9166 138 9200
rect 1572 9166 1588 9200
rect 122 9080 138 9114
rect 1572 9080 1588 9114
rect 122 8994 138 9028
rect 1572 8994 1588 9028
rect 122 8908 138 8942
rect 1572 8908 1588 8942
rect 122 8822 138 8856
rect 1572 8822 1588 8856
rect 122 8736 138 8770
rect 1572 8736 1588 8770
rect 122 8650 138 8684
rect 1572 8650 1588 8684
rect 122 8564 138 8598
rect 1572 8564 1588 8598
rect 122 8478 138 8512
rect 1572 8478 1588 8512
rect 122 8392 138 8426
rect 1572 8392 1588 8426
rect 122 8306 138 8340
rect 1572 8306 1588 8340
rect 122 8220 138 8254
rect 1572 8220 1588 8254
rect 122 8134 138 8168
rect 1572 8134 1588 8168
rect 122 8048 138 8082
rect 1572 8048 1588 8082
rect 122 7962 138 7996
rect 1572 7962 1588 7996
rect 122 7876 138 7910
rect 1572 7876 1588 7910
rect 122 7790 138 7824
rect 1572 7790 1588 7824
rect 122 7704 138 7738
rect 1572 7704 1588 7738
rect 122 7618 138 7652
rect 1572 7618 1588 7652
rect 122 7532 138 7566
rect 1572 7532 1588 7566
rect 122 7446 138 7480
rect 1572 7446 1588 7480
rect 122 7360 138 7394
rect 1572 7360 1588 7394
rect 122 7274 138 7308
rect 1572 7274 1588 7308
rect 122 7188 138 7222
rect 1572 7188 1588 7222
rect 122 7102 138 7136
rect 1572 7102 1588 7136
rect 122 7016 138 7050
rect 1572 7016 1588 7050
rect 122 6930 138 6964
rect 1572 6930 1588 6964
rect 122 6844 138 6878
rect 1572 6844 1588 6878
rect 122 6758 138 6792
rect 1572 6758 1588 6792
rect 122 6672 138 6706
rect 1572 6672 1588 6706
rect 122 6586 138 6620
rect 1572 6586 1588 6620
rect 122 6500 138 6534
rect 1572 6500 1588 6534
rect 122 6414 138 6448
rect 1572 6414 1588 6448
rect 122 6328 138 6362
rect 1572 6328 1588 6362
rect 122 6242 138 6276
rect 1572 6242 1588 6276
rect 122 6156 138 6190
rect 1572 6156 1588 6190
rect 122 6070 138 6104
rect 1572 6070 1588 6104
rect 122 5984 138 6018
rect 1572 5984 1588 6018
rect 122 5898 138 5932
rect 1572 5898 1588 5932
rect 122 5812 138 5846
rect 1572 5812 1588 5846
rect 122 5726 138 5760
rect 1572 5726 1588 5760
rect 122 5640 138 5674
rect 1572 5640 1588 5674
rect 122 5554 138 5588
rect 1572 5554 1588 5588
rect 122 5468 138 5502
rect 1572 5468 1588 5502
rect 122 5382 138 5416
rect 1572 5382 1588 5416
rect 122 5296 138 5330
rect 1572 5296 1588 5330
rect 122 5210 138 5244
rect 1572 5210 1588 5244
rect 122 5124 138 5158
rect 1572 5124 1588 5158
rect 122 5038 138 5072
rect 1572 5038 1588 5072
rect 122 4952 138 4986
rect 1572 4952 1588 4986
rect 122 4866 138 4900
rect 1572 4866 1588 4900
rect 122 4780 138 4814
rect 1572 4780 1588 4814
rect 122 4694 138 4728
rect 1572 4694 1588 4728
rect 122 4608 138 4642
rect 1572 4608 1588 4642
rect 122 4522 138 4556
rect 1572 4522 1588 4556
rect 122 4436 138 4470
rect 1572 4436 1588 4470
rect 122 4350 138 4384
rect 1572 4350 1588 4384
rect 122 4264 138 4298
rect 1572 4264 1588 4298
rect 122 4178 138 4212
rect 1572 4178 1588 4212
rect 122 4092 138 4126
rect 1572 4092 1588 4126
rect 122 4006 138 4040
rect 1572 4006 1588 4040
rect 122 3920 138 3954
rect 1572 3920 1588 3954
rect 122 3834 138 3868
rect 1572 3834 1588 3868
rect 122 3748 138 3782
rect 1572 3748 1588 3782
rect 122 3662 138 3696
rect 1572 3662 1588 3696
rect 122 3576 138 3610
rect 1572 3576 1588 3610
rect 122 3490 138 3524
rect 1572 3490 1588 3524
rect 122 3404 138 3438
rect 1572 3404 1588 3438
rect 122 3318 138 3352
rect 1572 3318 1588 3352
rect 122 3232 138 3266
rect 1572 3232 1588 3266
rect 122 3146 138 3180
rect 1572 3146 1588 3180
rect 122 3060 138 3094
rect 1572 3060 1588 3094
rect 122 2974 138 3008
rect 1572 2974 1588 3008
rect 122 2888 138 2922
rect 1572 2888 1588 2922
rect 122 2802 138 2836
rect 1572 2802 1588 2836
rect 122 2716 138 2750
rect 1572 2716 1588 2750
rect 122 2630 138 2664
rect 1572 2630 1588 2664
rect 122 2544 138 2578
rect 1572 2544 1588 2578
rect 122 2458 138 2492
rect 1572 2458 1588 2492
rect 122 2372 138 2406
rect 1572 2372 1588 2406
rect 122 2286 138 2320
rect 1572 2286 1588 2320
rect 122 2200 138 2234
rect 1572 2200 1588 2234
rect 122 2114 138 2148
rect 1572 2114 1588 2148
rect 122 2028 138 2062
rect 1572 2028 1588 2062
rect 122 1942 138 1976
rect 1572 1942 1588 1976
rect 122 1856 138 1890
rect 1572 1856 1588 1890
rect 122 1770 138 1804
rect 1572 1770 1588 1804
rect 122 1684 138 1718
rect 1572 1684 1588 1718
rect 122 1598 138 1632
rect 1572 1598 1588 1632
rect 122 1512 138 1546
rect 1572 1512 1588 1546
rect 122 1426 138 1460
rect 1572 1426 1588 1460
rect 122 1340 138 1374
rect 1572 1340 1588 1374
rect 122 1254 138 1288
rect 1572 1254 1588 1288
rect 122 1168 138 1202
rect 1572 1168 1588 1202
rect 122 1082 138 1116
rect 1572 1082 1588 1116
rect 122 996 138 1030
rect 1572 996 1588 1030
rect 122 910 138 944
rect 1572 910 1588 944
rect 122 824 138 858
rect 1572 824 1588 858
rect 122 738 138 772
rect 1572 738 1588 772
rect 122 652 138 686
rect 1572 652 1588 686
rect 122 566 138 600
rect 1572 566 1588 600
rect 122 480 138 514
rect 1572 480 1588 514
rect 122 394 138 428
rect 1572 394 1588 428
rect 122 308 138 342
rect 1572 308 1588 342
rect 122 222 138 256
rect 1572 222 1588 256
rect 122 136 138 170
rect 1572 136 1588 170
rect 1628 163 1662 179
rect 36 70 70 100
rect 1710 70 1744 100
rect 36 36 100 70
rect 1680 36 1744 70
<< viali >>
rect 100 100168 1680 100202
rect 36 100 70 100138
rect 138 100068 1572 100102
rect 138 99982 1572 100016
rect 138 99896 1572 99930
rect 138 99810 1572 99844
rect 138 99724 1572 99758
rect 138 99638 1572 99672
rect 138 99552 1572 99586
rect 138 99466 1572 99500
rect 138 99380 1572 99414
rect 138 99294 1572 99328
rect 138 99208 1572 99242
rect 138 99122 1572 99156
rect 138 99036 1572 99070
rect 138 98950 1572 98984
rect 138 98864 1572 98898
rect 138 98778 1572 98812
rect 138 98692 1572 98726
rect 138 98606 1572 98640
rect 138 98520 1572 98554
rect 138 98434 1572 98468
rect 138 98348 1572 98382
rect 138 98262 1572 98296
rect 138 98176 1572 98210
rect 138 98090 1572 98124
rect 138 98004 1572 98038
rect 138 97918 1572 97952
rect 138 97832 1572 97866
rect 138 97746 1572 97780
rect 138 97660 1572 97694
rect 138 97574 1572 97608
rect 138 97488 1572 97522
rect 138 97402 1572 97436
rect 138 97316 1572 97350
rect 138 97230 1572 97264
rect 138 97144 1572 97178
rect 138 97058 1572 97092
rect 138 96972 1572 97006
rect 138 96886 1572 96920
rect 138 96800 1572 96834
rect 138 96714 1572 96748
rect 138 96628 1572 96662
rect 138 96542 1572 96576
rect 138 96456 1572 96490
rect 138 96370 1572 96404
rect 138 96284 1572 96318
rect 138 96198 1572 96232
rect 138 96112 1572 96146
rect 138 96026 1572 96060
rect 138 95940 1572 95974
rect 138 95854 1572 95888
rect 138 95768 1572 95802
rect 138 95682 1572 95716
rect 138 95596 1572 95630
rect 138 95510 1572 95544
rect 138 95424 1572 95458
rect 138 95338 1572 95372
rect 138 95252 1572 95286
rect 138 95166 1572 95200
rect 138 95080 1572 95114
rect 138 94994 1572 95028
rect 138 94908 1572 94942
rect 138 94822 1572 94856
rect 138 94736 1572 94770
rect 138 94650 1572 94684
rect 138 94564 1572 94598
rect 138 94478 1572 94512
rect 138 94392 1572 94426
rect 138 94306 1572 94340
rect 138 94220 1572 94254
rect 138 94134 1572 94168
rect 138 94048 1572 94082
rect 138 93962 1572 93996
rect 138 93876 1572 93910
rect 138 93790 1572 93824
rect 138 93704 1572 93738
rect 138 93618 1572 93652
rect 138 93532 1572 93566
rect 138 93446 1572 93480
rect 138 93360 1572 93394
rect 138 93274 1572 93308
rect 138 93188 1572 93222
rect 138 93102 1572 93136
rect 138 93016 1572 93050
rect 138 92930 1572 92964
rect 138 92844 1572 92878
rect 138 92758 1572 92792
rect 138 92672 1572 92706
rect 138 92586 1572 92620
rect 138 92500 1572 92534
rect 138 92414 1572 92448
rect 138 92328 1572 92362
rect 138 92242 1572 92276
rect 138 92156 1572 92190
rect 138 92070 1572 92104
rect 138 91984 1572 92018
rect 138 91898 1572 91932
rect 138 91812 1572 91846
rect 138 91726 1572 91760
rect 138 91640 1572 91674
rect 138 91554 1572 91588
rect 138 91468 1572 91502
rect 138 91382 1572 91416
rect 138 91296 1572 91330
rect 138 91210 1572 91244
rect 138 91124 1572 91158
rect 138 91038 1572 91072
rect 138 90952 1572 90986
rect 138 90866 1572 90900
rect 138 90780 1572 90814
rect 138 90694 1572 90728
rect 138 90608 1572 90642
rect 138 90522 1572 90556
rect 138 90436 1572 90470
rect 138 90350 1572 90384
rect 138 90264 1572 90298
rect 138 90178 1572 90212
rect 138 90092 1572 90126
rect 138 90006 1572 90040
rect 138 89920 1572 89954
rect 138 89834 1572 89868
rect 138 89748 1572 89782
rect 138 89662 1572 89696
rect 138 89576 1572 89610
rect 138 89490 1572 89524
rect 138 89404 1572 89438
rect 138 89318 1572 89352
rect 138 89232 1572 89266
rect 138 89146 1572 89180
rect 138 89060 1572 89094
rect 138 88974 1572 89008
rect 138 88888 1572 88922
rect 138 88802 1572 88836
rect 138 88716 1572 88750
rect 138 88630 1572 88664
rect 138 88544 1572 88578
rect 138 88458 1572 88492
rect 138 88372 1572 88406
rect 138 88286 1572 88320
rect 138 88200 1572 88234
rect 138 88114 1572 88148
rect 138 88028 1572 88062
rect 138 87942 1572 87976
rect 138 87856 1572 87890
rect 138 87770 1572 87804
rect 138 87684 1572 87718
rect 138 87598 1572 87632
rect 138 87512 1572 87546
rect 138 87426 1572 87460
rect 138 87340 1572 87374
rect 138 87254 1572 87288
rect 138 87168 1572 87202
rect 138 87082 1572 87116
rect 138 86996 1572 87030
rect 138 86910 1572 86944
rect 138 86824 1572 86858
rect 138 86738 1572 86772
rect 138 86652 1572 86686
rect 138 86566 1572 86600
rect 138 86480 1572 86514
rect 138 86394 1572 86428
rect 138 86308 1572 86342
rect 138 86222 1572 86256
rect 138 86136 1572 86170
rect 138 86050 1572 86084
rect 138 85964 1572 85998
rect 138 85878 1572 85912
rect 138 85792 1572 85826
rect 138 85706 1572 85740
rect 138 85620 1572 85654
rect 138 85534 1572 85568
rect 138 85448 1572 85482
rect 138 85362 1572 85396
rect 138 85276 1572 85310
rect 138 85190 1572 85224
rect 138 85104 1572 85138
rect 138 85018 1572 85052
rect 138 84932 1572 84966
rect 138 84846 1572 84880
rect 138 84760 1572 84794
rect 138 84674 1572 84708
rect 138 84588 1572 84622
rect 138 84502 1572 84536
rect 138 84416 1572 84450
rect 138 84330 1572 84364
rect 138 84244 1572 84278
rect 138 84158 1572 84192
rect 138 84072 1572 84106
rect 138 83986 1572 84020
rect 138 83900 1572 83934
rect 138 83814 1572 83848
rect 138 83728 1572 83762
rect 138 83642 1572 83676
rect 138 83556 1572 83590
rect 138 83470 1572 83504
rect 138 83384 1572 83418
rect 138 83298 1572 83332
rect 138 83212 1572 83246
rect 138 83126 1572 83160
rect 138 83040 1572 83074
rect 138 82954 1572 82988
rect 138 82868 1572 82902
rect 138 82782 1572 82816
rect 138 82696 1572 82730
rect 138 82610 1572 82644
rect 138 82524 1572 82558
rect 138 82438 1572 82472
rect 138 82352 1572 82386
rect 138 82266 1572 82300
rect 138 82180 1572 82214
rect 138 82094 1572 82128
rect 138 82008 1572 82042
rect 138 81922 1572 81956
rect 138 81836 1572 81870
rect 138 81750 1572 81784
rect 138 81664 1572 81698
rect 138 81578 1572 81612
rect 138 81492 1572 81526
rect 138 81406 1572 81440
rect 138 81320 1572 81354
rect 138 81234 1572 81268
rect 138 81148 1572 81182
rect 138 81062 1572 81096
rect 138 80976 1572 81010
rect 138 80890 1572 80924
rect 138 80804 1572 80838
rect 138 80718 1572 80752
rect 138 80632 1572 80666
rect 138 80546 1572 80580
rect 138 80460 1572 80494
rect 138 80374 1572 80408
rect 138 80288 1572 80322
rect 138 80202 1572 80236
rect 138 80116 1572 80150
rect 138 80030 1572 80064
rect 138 79944 1572 79978
rect 138 79858 1572 79892
rect 138 79772 1572 79806
rect 138 79686 1572 79720
rect 138 79600 1572 79634
rect 138 79514 1572 79548
rect 138 79428 1572 79462
rect 138 79342 1572 79376
rect 138 79256 1572 79290
rect 138 79170 1572 79204
rect 138 79084 1572 79118
rect 138 78998 1572 79032
rect 138 78912 1572 78946
rect 138 78826 1572 78860
rect 138 78740 1572 78774
rect 138 78654 1572 78688
rect 138 78568 1572 78602
rect 138 78482 1572 78516
rect 138 78396 1572 78430
rect 138 78310 1572 78344
rect 138 78224 1572 78258
rect 138 78138 1572 78172
rect 138 78052 1572 78086
rect 138 77966 1572 78000
rect 138 77880 1572 77914
rect 138 77794 1572 77828
rect 138 77708 1572 77742
rect 138 77622 1572 77656
rect 138 77536 1572 77570
rect 138 77450 1572 77484
rect 138 77364 1572 77398
rect 138 77278 1572 77312
rect 138 77192 1572 77226
rect 138 77106 1572 77140
rect 138 77020 1572 77054
rect 138 76934 1572 76968
rect 138 76848 1572 76882
rect 138 76762 1572 76796
rect 138 76676 1572 76710
rect 138 76590 1572 76624
rect 138 76504 1572 76538
rect 138 76418 1572 76452
rect 138 76332 1572 76366
rect 138 76246 1572 76280
rect 138 76160 1572 76194
rect 138 76074 1572 76108
rect 138 75988 1572 76022
rect 138 75902 1572 75936
rect 138 75816 1572 75850
rect 138 75730 1572 75764
rect 138 75644 1572 75678
rect 138 75558 1572 75592
rect 138 75472 1572 75506
rect 138 75386 1572 75420
rect 138 75300 1572 75334
rect 138 75214 1572 75248
rect 138 75128 1572 75162
rect 138 75042 1572 75076
rect 138 74956 1572 74990
rect 138 74870 1572 74904
rect 138 74784 1572 74818
rect 138 74698 1572 74732
rect 138 74612 1572 74646
rect 138 74526 1572 74560
rect 138 74440 1572 74474
rect 138 74354 1572 74388
rect 138 74268 1572 74302
rect 138 74182 1572 74216
rect 138 74096 1572 74130
rect 138 74010 1572 74044
rect 138 73924 1572 73958
rect 138 73838 1572 73872
rect 138 73752 1572 73786
rect 138 73666 1572 73700
rect 138 73580 1572 73614
rect 138 73494 1572 73528
rect 138 73408 1572 73442
rect 138 73322 1572 73356
rect 138 73236 1572 73270
rect 138 73150 1572 73184
rect 138 73064 1572 73098
rect 138 72978 1572 73012
rect 138 72892 1572 72926
rect 138 72806 1572 72840
rect 138 72720 1572 72754
rect 138 72634 1572 72668
rect 138 72548 1572 72582
rect 138 72462 1572 72496
rect 138 72376 1572 72410
rect 138 72290 1572 72324
rect 138 72204 1572 72238
rect 138 72118 1572 72152
rect 138 72032 1572 72066
rect 138 71946 1572 71980
rect 138 71860 1572 71894
rect 138 71774 1572 71808
rect 138 71688 1572 71722
rect 138 71602 1572 71636
rect 138 71516 1572 71550
rect 138 71430 1572 71464
rect 138 71344 1572 71378
rect 138 71258 1572 71292
rect 138 71172 1572 71206
rect 138 71086 1572 71120
rect 138 71000 1572 71034
rect 138 70914 1572 70948
rect 138 70828 1572 70862
rect 138 70742 1572 70776
rect 138 70656 1572 70690
rect 138 70570 1572 70604
rect 138 70484 1572 70518
rect 138 70398 1572 70432
rect 138 70312 1572 70346
rect 138 70226 1572 70260
rect 138 70140 1572 70174
rect 138 70054 1572 70088
rect 138 69968 1572 70002
rect 138 69882 1572 69916
rect 138 69796 1572 69830
rect 138 69710 1572 69744
rect 138 69624 1572 69658
rect 138 69538 1572 69572
rect 138 69452 1572 69486
rect 138 69366 1572 69400
rect 138 69280 1572 69314
rect 138 69194 1572 69228
rect 138 69108 1572 69142
rect 138 69022 1572 69056
rect 138 68936 1572 68970
rect 138 68850 1572 68884
rect 138 68764 1572 68798
rect 138 68678 1572 68712
rect 138 68592 1572 68626
rect 138 68506 1572 68540
rect 138 68420 1572 68454
rect 138 68334 1572 68368
rect 138 68248 1572 68282
rect 138 68162 1572 68196
rect 138 68076 1572 68110
rect 138 67990 1572 68024
rect 138 67904 1572 67938
rect 138 67818 1572 67852
rect 138 67732 1572 67766
rect 138 67646 1572 67680
rect 138 67560 1572 67594
rect 138 67474 1572 67508
rect 138 67388 1572 67422
rect 138 67302 1572 67336
rect 138 67216 1572 67250
rect 138 67130 1572 67164
rect 138 67044 1572 67078
rect 138 66958 1572 66992
rect 138 66872 1572 66906
rect 138 66786 1572 66820
rect 138 66700 1572 66734
rect 138 66614 1572 66648
rect 138 66528 1572 66562
rect 138 66442 1572 66476
rect 138 66356 1572 66390
rect 138 66270 1572 66304
rect 138 66184 1572 66218
rect 138 66098 1572 66132
rect 138 66012 1572 66046
rect 138 65926 1572 65960
rect 138 65840 1572 65874
rect 138 65754 1572 65788
rect 138 65668 1572 65702
rect 138 65582 1572 65616
rect 138 65496 1572 65530
rect 138 65410 1572 65444
rect 138 65324 1572 65358
rect 138 65238 1572 65272
rect 138 65152 1572 65186
rect 138 65066 1572 65100
rect 138 64980 1572 65014
rect 138 64894 1572 64928
rect 138 64808 1572 64842
rect 138 64722 1572 64756
rect 138 64636 1572 64670
rect 138 64550 1572 64584
rect 138 64464 1572 64498
rect 138 64378 1572 64412
rect 138 64292 1572 64326
rect 138 64206 1572 64240
rect 138 64120 1572 64154
rect 138 64034 1572 64068
rect 138 63948 1572 63982
rect 138 63862 1572 63896
rect 138 63776 1572 63810
rect 138 63690 1572 63724
rect 138 63604 1572 63638
rect 138 63518 1572 63552
rect 138 63432 1572 63466
rect 138 63346 1572 63380
rect 138 63260 1572 63294
rect 138 63174 1572 63208
rect 138 63088 1572 63122
rect 138 63002 1572 63036
rect 138 62916 1572 62950
rect 138 62830 1572 62864
rect 138 62744 1572 62778
rect 138 62658 1572 62692
rect 138 62572 1572 62606
rect 138 62486 1572 62520
rect 138 62400 1572 62434
rect 138 62314 1572 62348
rect 138 62228 1572 62262
rect 138 62142 1572 62176
rect 138 62056 1572 62090
rect 138 61970 1572 62004
rect 138 61884 1572 61918
rect 138 61798 1572 61832
rect 138 61712 1572 61746
rect 138 61626 1572 61660
rect 138 61540 1572 61574
rect 138 61454 1572 61488
rect 138 61368 1572 61402
rect 138 61282 1572 61316
rect 138 61196 1572 61230
rect 138 61110 1572 61144
rect 138 61024 1572 61058
rect 138 60938 1572 60972
rect 138 60852 1572 60886
rect 138 60766 1572 60800
rect 138 60680 1572 60714
rect 138 60594 1572 60628
rect 138 60508 1572 60542
rect 138 60422 1572 60456
rect 138 60336 1572 60370
rect 138 60250 1572 60284
rect 138 60164 1572 60198
rect 138 60078 1572 60112
rect 138 59992 1572 60026
rect 138 59906 1572 59940
rect 138 59820 1572 59854
rect 138 59734 1572 59768
rect 138 59648 1572 59682
rect 138 59562 1572 59596
rect 138 59476 1572 59510
rect 138 59390 1572 59424
rect 138 59304 1572 59338
rect 138 59218 1572 59252
rect 138 59132 1572 59166
rect 138 59046 1572 59080
rect 138 58960 1572 58994
rect 138 58874 1572 58908
rect 138 58788 1572 58822
rect 138 58702 1572 58736
rect 138 58616 1572 58650
rect 138 58530 1572 58564
rect 138 58444 1572 58478
rect 138 58358 1572 58392
rect 138 58272 1572 58306
rect 138 58186 1572 58220
rect 138 58100 1572 58134
rect 138 58014 1572 58048
rect 138 57928 1572 57962
rect 138 57842 1572 57876
rect 138 57756 1572 57790
rect 138 57670 1572 57704
rect 138 57584 1572 57618
rect 138 57498 1572 57532
rect 138 57412 1572 57446
rect 138 57326 1572 57360
rect 138 57240 1572 57274
rect 138 57154 1572 57188
rect 138 57068 1572 57102
rect 138 56982 1572 57016
rect 138 56896 1572 56930
rect 138 56810 1572 56844
rect 138 56724 1572 56758
rect 138 56638 1572 56672
rect 138 56552 1572 56586
rect 138 56466 1572 56500
rect 138 56380 1572 56414
rect 138 56294 1572 56328
rect 138 56208 1572 56242
rect 138 56122 1572 56156
rect 138 56036 1572 56070
rect 138 55950 1572 55984
rect 138 55864 1572 55898
rect 138 55778 1572 55812
rect 138 55692 1572 55726
rect 138 55606 1572 55640
rect 138 55520 1572 55554
rect 138 55434 1572 55468
rect 138 55348 1572 55382
rect 138 55262 1572 55296
rect 138 55176 1572 55210
rect 138 55090 1572 55124
rect 138 55004 1572 55038
rect 138 54918 1572 54952
rect 138 54832 1572 54866
rect 138 54746 1572 54780
rect 138 54660 1572 54694
rect 138 54574 1572 54608
rect 138 54488 1572 54522
rect 138 54402 1572 54436
rect 138 54316 1572 54350
rect 138 54230 1572 54264
rect 138 54144 1572 54178
rect 138 54058 1572 54092
rect 138 53972 1572 54006
rect 138 53886 1572 53920
rect 138 53800 1572 53834
rect 138 53714 1572 53748
rect 138 53628 1572 53662
rect 138 53542 1572 53576
rect 138 53456 1572 53490
rect 138 53370 1572 53404
rect 138 53284 1572 53318
rect 138 53198 1572 53232
rect 138 53112 1572 53146
rect 138 53026 1572 53060
rect 138 52940 1572 52974
rect 138 52854 1572 52888
rect 138 52768 1572 52802
rect 138 52682 1572 52716
rect 138 52596 1572 52630
rect 138 52510 1572 52544
rect 138 52424 1572 52458
rect 138 52338 1572 52372
rect 138 52252 1572 52286
rect 138 52166 1572 52200
rect 138 52080 1572 52114
rect 138 51994 1572 52028
rect 138 51908 1572 51942
rect 138 51822 1572 51856
rect 138 51736 1572 51770
rect 138 51650 1572 51684
rect 138 51564 1572 51598
rect 138 51478 1572 51512
rect 138 51392 1572 51426
rect 138 51306 1572 51340
rect 138 51220 1572 51254
rect 138 51134 1572 51168
rect 138 51048 1572 51082
rect 138 50962 1572 50996
rect 138 50876 1572 50910
rect 138 50790 1572 50824
rect 138 50704 1572 50738
rect 138 50618 1572 50652
rect 138 50532 1572 50566
rect 138 50446 1572 50480
rect 138 50360 1572 50394
rect 138 50274 1572 50308
rect 138 50188 1572 50222
rect 138 50102 1572 50136
rect 138 50016 1572 50050
rect 138 49930 1572 49964
rect 138 49844 1572 49878
rect 138 49758 1572 49792
rect 138 49672 1572 49706
rect 138 49586 1572 49620
rect 138 49500 1572 49534
rect 138 49414 1572 49448
rect 138 49328 1572 49362
rect 138 49242 1572 49276
rect 138 49156 1572 49190
rect 138 49070 1572 49104
rect 138 48984 1572 49018
rect 138 48898 1572 48932
rect 138 48812 1572 48846
rect 138 48726 1572 48760
rect 138 48640 1572 48674
rect 138 48554 1572 48588
rect 138 48468 1572 48502
rect 138 48382 1572 48416
rect 138 48296 1572 48330
rect 138 48210 1572 48244
rect 138 48124 1572 48158
rect 138 48038 1572 48072
rect 138 47952 1572 47986
rect 138 47866 1572 47900
rect 138 47780 1572 47814
rect 138 47694 1572 47728
rect 138 47608 1572 47642
rect 138 47522 1572 47556
rect 138 47436 1572 47470
rect 138 47350 1572 47384
rect 138 47264 1572 47298
rect 138 47178 1572 47212
rect 138 47092 1572 47126
rect 138 47006 1572 47040
rect 138 46920 1572 46954
rect 138 46834 1572 46868
rect 138 46748 1572 46782
rect 138 46662 1572 46696
rect 138 46576 1572 46610
rect 138 46490 1572 46524
rect 138 46404 1572 46438
rect 138 46318 1572 46352
rect 138 46232 1572 46266
rect 138 46146 1572 46180
rect 138 46060 1572 46094
rect 138 45974 1572 46008
rect 138 45888 1572 45922
rect 138 45802 1572 45836
rect 138 45716 1572 45750
rect 138 45630 1572 45664
rect 138 45544 1572 45578
rect 138 45458 1572 45492
rect 138 45372 1572 45406
rect 138 45286 1572 45320
rect 138 45200 1572 45234
rect 138 45114 1572 45148
rect 138 45028 1572 45062
rect 138 44942 1572 44976
rect 138 44856 1572 44890
rect 138 44770 1572 44804
rect 138 44684 1572 44718
rect 138 44598 1572 44632
rect 138 44512 1572 44546
rect 138 44426 1572 44460
rect 138 44340 1572 44374
rect 138 44254 1572 44288
rect 138 44168 1572 44202
rect 138 44082 1572 44116
rect 138 43996 1572 44030
rect 138 43910 1572 43944
rect 138 43824 1572 43858
rect 138 43738 1572 43772
rect 138 43652 1572 43686
rect 138 43566 1572 43600
rect 138 43480 1572 43514
rect 138 43394 1572 43428
rect 138 43308 1572 43342
rect 138 43222 1572 43256
rect 138 43136 1572 43170
rect 138 43050 1572 43084
rect 138 42964 1572 42998
rect 138 42878 1572 42912
rect 138 42792 1572 42826
rect 138 42706 1572 42740
rect 138 42620 1572 42654
rect 138 42534 1572 42568
rect 138 42448 1572 42482
rect 138 42362 1572 42396
rect 138 42276 1572 42310
rect 138 42190 1572 42224
rect 138 42104 1572 42138
rect 138 42018 1572 42052
rect 138 41932 1572 41966
rect 138 41846 1572 41880
rect 138 41760 1572 41794
rect 138 41674 1572 41708
rect 138 41588 1572 41622
rect 138 41502 1572 41536
rect 138 41416 1572 41450
rect 138 41330 1572 41364
rect 138 41244 1572 41278
rect 138 41158 1572 41192
rect 138 41072 1572 41106
rect 138 40986 1572 41020
rect 138 40900 1572 40934
rect 138 40814 1572 40848
rect 138 40728 1572 40762
rect 138 40642 1572 40676
rect 138 40556 1572 40590
rect 138 40470 1572 40504
rect 138 40384 1572 40418
rect 138 40298 1572 40332
rect 138 40212 1572 40246
rect 138 40126 1572 40160
rect 138 40040 1572 40074
rect 138 39954 1572 39988
rect 138 39868 1572 39902
rect 138 39782 1572 39816
rect 138 39696 1572 39730
rect 138 39610 1572 39644
rect 138 39524 1572 39558
rect 138 39438 1572 39472
rect 138 39352 1572 39386
rect 138 39266 1572 39300
rect 138 39180 1572 39214
rect 138 39094 1572 39128
rect 138 39008 1572 39042
rect 138 38922 1572 38956
rect 138 38836 1572 38870
rect 138 38750 1572 38784
rect 138 38664 1572 38698
rect 138 38578 1572 38612
rect 138 38492 1572 38526
rect 138 38406 1572 38440
rect 138 38320 1572 38354
rect 138 38234 1572 38268
rect 138 38148 1572 38182
rect 138 38062 1572 38096
rect 138 37976 1572 38010
rect 138 37890 1572 37924
rect 138 37804 1572 37838
rect 138 37718 1572 37752
rect 138 37632 1572 37666
rect 138 37546 1572 37580
rect 138 37460 1572 37494
rect 138 37374 1572 37408
rect 138 37288 1572 37322
rect 138 37202 1572 37236
rect 138 37116 1572 37150
rect 138 37030 1572 37064
rect 138 36944 1572 36978
rect 138 36858 1572 36892
rect 138 36772 1572 36806
rect 138 36686 1572 36720
rect 138 36600 1572 36634
rect 138 36514 1572 36548
rect 138 36428 1572 36462
rect 138 36342 1572 36376
rect 138 36256 1572 36290
rect 138 36170 1572 36204
rect 138 36084 1572 36118
rect 138 35998 1572 36032
rect 138 35912 1572 35946
rect 138 35826 1572 35860
rect 138 35740 1572 35774
rect 138 35654 1572 35688
rect 138 35568 1572 35602
rect 138 35482 1572 35516
rect 138 35396 1572 35430
rect 138 35310 1572 35344
rect 138 35224 1572 35258
rect 138 35138 1572 35172
rect 138 35052 1572 35086
rect 138 34966 1572 35000
rect 138 34880 1572 34914
rect 138 34794 1572 34828
rect 138 34708 1572 34742
rect 138 34622 1572 34656
rect 138 34536 1572 34570
rect 138 34450 1572 34484
rect 138 34364 1572 34398
rect 138 34278 1572 34312
rect 138 34192 1572 34226
rect 138 34106 1572 34140
rect 138 34020 1572 34054
rect 138 33934 1572 33968
rect 138 33848 1572 33882
rect 138 33762 1572 33796
rect 138 33676 1572 33710
rect 138 33590 1572 33624
rect 138 33504 1572 33538
rect 138 33418 1572 33452
rect 138 33332 1572 33366
rect 138 33246 1572 33280
rect 138 33160 1572 33194
rect 138 33074 1572 33108
rect 138 32988 1572 33022
rect 138 32902 1572 32936
rect 138 32816 1572 32850
rect 138 32730 1572 32764
rect 138 32644 1572 32678
rect 138 32558 1572 32592
rect 138 32472 1572 32506
rect 138 32386 1572 32420
rect 138 32300 1572 32334
rect 138 32214 1572 32248
rect 138 32128 1572 32162
rect 138 32042 1572 32076
rect 138 31956 1572 31990
rect 138 31870 1572 31904
rect 138 31784 1572 31818
rect 138 31698 1572 31732
rect 138 31612 1572 31646
rect 138 31526 1572 31560
rect 138 31440 1572 31474
rect 138 31354 1572 31388
rect 138 31268 1572 31302
rect 138 31182 1572 31216
rect 138 31096 1572 31130
rect 138 31010 1572 31044
rect 138 30924 1572 30958
rect 138 30838 1572 30872
rect 138 30752 1572 30786
rect 138 30666 1572 30700
rect 138 30580 1572 30614
rect 138 30494 1572 30528
rect 138 30408 1572 30442
rect 138 30322 1572 30356
rect 138 30236 1572 30270
rect 138 30150 1572 30184
rect 138 30064 1572 30098
rect 138 29978 1572 30012
rect 138 29892 1572 29926
rect 138 29806 1572 29840
rect 138 29720 1572 29754
rect 138 29634 1572 29668
rect 138 29548 1572 29582
rect 138 29462 1572 29496
rect 138 29376 1572 29410
rect 138 29290 1572 29324
rect 138 29204 1572 29238
rect 138 29118 1572 29152
rect 138 29032 1572 29066
rect 138 28946 1572 28980
rect 138 28860 1572 28894
rect 138 28774 1572 28808
rect 138 28688 1572 28722
rect 138 28602 1572 28636
rect 138 28516 1572 28550
rect 138 28430 1572 28464
rect 138 28344 1572 28378
rect 138 28258 1572 28292
rect 138 28172 1572 28206
rect 138 28086 1572 28120
rect 138 28000 1572 28034
rect 138 27914 1572 27948
rect 138 27828 1572 27862
rect 138 27742 1572 27776
rect 138 27656 1572 27690
rect 138 27570 1572 27604
rect 138 27484 1572 27518
rect 138 27398 1572 27432
rect 138 27312 1572 27346
rect 138 27226 1572 27260
rect 138 27140 1572 27174
rect 138 27054 1572 27088
rect 138 26968 1572 27002
rect 138 26882 1572 26916
rect 138 26796 1572 26830
rect 138 26710 1572 26744
rect 138 26624 1572 26658
rect 138 26538 1572 26572
rect 138 26452 1572 26486
rect 138 26366 1572 26400
rect 138 26280 1572 26314
rect 138 26194 1572 26228
rect 138 26108 1572 26142
rect 138 26022 1572 26056
rect 138 25936 1572 25970
rect 138 25850 1572 25884
rect 138 25764 1572 25798
rect 138 25678 1572 25712
rect 138 25592 1572 25626
rect 138 25506 1572 25540
rect 138 25420 1572 25454
rect 138 25334 1572 25368
rect 138 25248 1572 25282
rect 138 25162 1572 25196
rect 138 25076 1572 25110
rect 138 24990 1572 25024
rect 138 24904 1572 24938
rect 138 24818 1572 24852
rect 138 24732 1572 24766
rect 138 24646 1572 24680
rect 138 24560 1572 24594
rect 138 24474 1572 24508
rect 138 24388 1572 24422
rect 138 24302 1572 24336
rect 138 24216 1572 24250
rect 138 24130 1572 24164
rect 138 24044 1572 24078
rect 138 23958 1572 23992
rect 138 23872 1572 23906
rect 138 23786 1572 23820
rect 138 23700 1572 23734
rect 138 23614 1572 23648
rect 138 23528 1572 23562
rect 138 23442 1572 23476
rect 138 23356 1572 23390
rect 138 23270 1572 23304
rect 138 23184 1572 23218
rect 138 23098 1572 23132
rect 138 23012 1572 23046
rect 138 22926 1572 22960
rect 138 22840 1572 22874
rect 138 22754 1572 22788
rect 138 22668 1572 22702
rect 138 22582 1572 22616
rect 138 22496 1572 22530
rect 138 22410 1572 22444
rect 138 22324 1572 22358
rect 138 22238 1572 22272
rect 138 22152 1572 22186
rect 138 22066 1572 22100
rect 138 21980 1572 22014
rect 138 21894 1572 21928
rect 138 21808 1572 21842
rect 138 21722 1572 21756
rect 138 21636 1572 21670
rect 138 21550 1572 21584
rect 138 21464 1572 21498
rect 138 21378 1572 21412
rect 138 21292 1572 21326
rect 138 21206 1572 21240
rect 138 21120 1572 21154
rect 138 21034 1572 21068
rect 138 20948 1572 20982
rect 138 20862 1572 20896
rect 138 20776 1572 20810
rect 138 20690 1572 20724
rect 138 20604 1572 20638
rect 138 20518 1572 20552
rect 138 20432 1572 20466
rect 138 20346 1572 20380
rect 138 20260 1572 20294
rect 138 20174 1572 20208
rect 138 20088 1572 20122
rect 138 20002 1572 20036
rect 138 19916 1572 19950
rect 138 19830 1572 19864
rect 138 19744 1572 19778
rect 138 19658 1572 19692
rect 138 19572 1572 19606
rect 138 19486 1572 19520
rect 138 19400 1572 19434
rect 138 19314 1572 19348
rect 138 19228 1572 19262
rect 138 19142 1572 19176
rect 138 19056 1572 19090
rect 138 18970 1572 19004
rect 138 18884 1572 18918
rect 138 18798 1572 18832
rect 138 18712 1572 18746
rect 138 18626 1572 18660
rect 138 18540 1572 18574
rect 138 18454 1572 18488
rect 138 18368 1572 18402
rect 138 18282 1572 18316
rect 138 18196 1572 18230
rect 138 18110 1572 18144
rect 138 18024 1572 18058
rect 138 17938 1572 17972
rect 138 17852 1572 17886
rect 138 17766 1572 17800
rect 138 17680 1572 17714
rect 138 17594 1572 17628
rect 138 17508 1572 17542
rect 138 17422 1572 17456
rect 138 17336 1572 17370
rect 138 17250 1572 17284
rect 138 17164 1572 17198
rect 138 17078 1572 17112
rect 138 16992 1572 17026
rect 138 16906 1572 16940
rect 138 16820 1572 16854
rect 138 16734 1572 16768
rect 138 16648 1572 16682
rect 138 16562 1572 16596
rect 138 16476 1572 16510
rect 138 16390 1572 16424
rect 138 16304 1572 16338
rect 138 16218 1572 16252
rect 138 16132 1572 16166
rect 138 16046 1572 16080
rect 138 15960 1572 15994
rect 138 15874 1572 15908
rect 138 15788 1572 15822
rect 138 15702 1572 15736
rect 138 15616 1572 15650
rect 138 15530 1572 15564
rect 138 15444 1572 15478
rect 138 15358 1572 15392
rect 138 15272 1572 15306
rect 138 15186 1572 15220
rect 138 15100 1572 15134
rect 138 15014 1572 15048
rect 138 14928 1572 14962
rect 138 14842 1572 14876
rect 138 14756 1572 14790
rect 138 14670 1572 14704
rect 138 14584 1572 14618
rect 138 14498 1572 14532
rect 138 14412 1572 14446
rect 138 14326 1572 14360
rect 138 14240 1572 14274
rect 138 14154 1572 14188
rect 138 14068 1572 14102
rect 138 13982 1572 14016
rect 138 13896 1572 13930
rect 138 13810 1572 13844
rect 138 13724 1572 13758
rect 138 13638 1572 13672
rect 138 13552 1572 13586
rect 138 13466 1572 13500
rect 138 13380 1572 13414
rect 138 13294 1572 13328
rect 138 13208 1572 13242
rect 138 13122 1572 13156
rect 138 13036 1572 13070
rect 138 12950 1572 12984
rect 138 12864 1572 12898
rect 138 12778 1572 12812
rect 138 12692 1572 12726
rect 138 12606 1572 12640
rect 138 12520 1572 12554
rect 138 12434 1572 12468
rect 138 12348 1572 12382
rect 138 12262 1572 12296
rect 138 12176 1572 12210
rect 138 12090 1572 12124
rect 138 12004 1572 12038
rect 138 11918 1572 11952
rect 138 11832 1572 11866
rect 138 11746 1572 11780
rect 138 11660 1572 11694
rect 138 11574 1572 11608
rect 138 11488 1572 11522
rect 138 11402 1572 11436
rect 138 11316 1572 11350
rect 138 11230 1572 11264
rect 138 11144 1572 11178
rect 138 11058 1572 11092
rect 138 10972 1572 11006
rect 138 10886 1572 10920
rect 138 10800 1572 10834
rect 138 10714 1572 10748
rect 138 10628 1572 10662
rect 138 10542 1572 10576
rect 138 10456 1572 10490
rect 138 10370 1572 10404
rect 138 10284 1572 10318
rect 138 10198 1572 10232
rect 138 10112 1572 10146
rect 138 10026 1572 10060
rect 138 9940 1572 9974
rect 138 9854 1572 9888
rect 138 9768 1572 9802
rect 138 9682 1572 9716
rect 138 9596 1572 9630
rect 138 9510 1572 9544
rect 138 9424 1572 9458
rect 138 9338 1572 9372
rect 138 9252 1572 9286
rect 138 9166 1572 9200
rect 138 9080 1572 9114
rect 138 8994 1572 9028
rect 138 8908 1572 8942
rect 138 8822 1572 8856
rect 138 8736 1572 8770
rect 138 8650 1572 8684
rect 138 8564 1572 8598
rect 138 8478 1572 8512
rect 138 8392 1572 8426
rect 138 8306 1572 8340
rect 138 8220 1572 8254
rect 138 8134 1572 8168
rect 138 8048 1572 8082
rect 138 7962 1572 7996
rect 138 7876 1572 7910
rect 138 7790 1572 7824
rect 138 7704 1572 7738
rect 138 7618 1572 7652
rect 138 7532 1572 7566
rect 138 7446 1572 7480
rect 138 7360 1572 7394
rect 138 7274 1572 7308
rect 138 7188 1572 7222
rect 138 7102 1572 7136
rect 138 7016 1572 7050
rect 138 6930 1572 6964
rect 138 6844 1572 6878
rect 138 6758 1572 6792
rect 138 6672 1572 6706
rect 138 6586 1572 6620
rect 138 6500 1572 6534
rect 138 6414 1572 6448
rect 138 6328 1572 6362
rect 138 6242 1572 6276
rect 138 6156 1572 6190
rect 138 6070 1572 6104
rect 138 5984 1572 6018
rect 138 5898 1572 5932
rect 138 5812 1572 5846
rect 138 5726 1572 5760
rect 138 5640 1572 5674
rect 138 5554 1572 5588
rect 138 5468 1572 5502
rect 138 5382 1572 5416
rect 138 5296 1572 5330
rect 138 5210 1572 5244
rect 138 5124 1572 5158
rect 138 5038 1572 5072
rect 138 4952 1572 4986
rect 138 4866 1572 4900
rect 138 4780 1572 4814
rect 138 4694 1572 4728
rect 138 4608 1572 4642
rect 138 4522 1572 4556
rect 138 4436 1572 4470
rect 138 4350 1572 4384
rect 138 4264 1572 4298
rect 138 4178 1572 4212
rect 138 4092 1572 4126
rect 138 4006 1572 4040
rect 138 3920 1572 3954
rect 138 3834 1572 3868
rect 138 3748 1572 3782
rect 138 3662 1572 3696
rect 138 3576 1572 3610
rect 138 3490 1572 3524
rect 138 3404 1572 3438
rect 138 3318 1572 3352
rect 138 3232 1572 3266
rect 138 3146 1572 3180
rect 138 3060 1572 3094
rect 138 2974 1572 3008
rect 138 2888 1572 2922
rect 138 2802 1572 2836
rect 138 2716 1572 2750
rect 138 2630 1572 2664
rect 138 2544 1572 2578
rect 138 2458 1572 2492
rect 138 2372 1572 2406
rect 138 2286 1572 2320
rect 138 2200 1572 2234
rect 138 2114 1572 2148
rect 138 2028 1572 2062
rect 138 1942 1572 1976
rect 138 1856 1572 1890
rect 138 1770 1572 1804
rect 138 1684 1572 1718
rect 138 1598 1572 1632
rect 138 1512 1572 1546
rect 138 1426 1572 1460
rect 138 1340 1572 1374
rect 138 1254 1572 1288
rect 138 1168 1572 1202
rect 138 1082 1572 1116
rect 138 996 1572 1030
rect 138 910 1572 944
rect 138 824 1572 858
rect 138 738 1572 772
rect 138 652 1572 686
rect 138 566 1572 600
rect 138 480 1572 514
rect 138 394 1572 428
rect 138 308 1572 342
rect 138 222 1572 256
rect 1628 179 1662 100059
rect 138 136 1572 170
rect 1710 100 1744 100138
rect 100 36 1680 70
<< metal1 >>
rect 30 100202 1750 100208
rect 30 100168 100 100202
rect 1680 100168 1750 100202
rect 30 100162 1750 100168
rect 30 100138 76 100162
rect 30 100 36 100138
rect 70 100 76 100138
rect 1704 100138 1750 100162
rect 894 100108 900 100111
rect 126 100102 900 100108
rect 1548 100108 1554 100111
rect 1548 100102 1584 100108
rect 126 100068 138 100102
rect 1572 100068 1584 100102
rect 126 100062 900 100068
rect 894 100059 900 100062
rect 1548 100062 1584 100068
rect 1618 100069 1672 100075
rect 1548 100059 1554 100062
rect 156 100022 162 100025
rect 126 100016 162 100022
rect 810 100022 816 100025
rect 810 100016 1584 100022
rect 126 99982 138 100016
rect 1572 99982 1584 100016
rect 126 99976 162 99982
rect 156 99973 162 99976
rect 810 99976 1584 99982
rect 810 99973 816 99976
rect 894 99936 900 99939
rect 126 99930 900 99936
rect 1548 99936 1554 99939
rect 1548 99930 1584 99936
rect 126 99896 138 99930
rect 1572 99896 1584 99930
rect 126 99890 900 99896
rect 894 99887 900 99890
rect 1548 99890 1584 99896
rect 1548 99887 1554 99890
rect 156 99850 162 99853
rect 126 99844 162 99850
rect 810 99850 816 99853
rect 810 99844 1584 99850
rect 126 99810 138 99844
rect 1572 99810 1584 99844
rect 126 99804 162 99810
rect 156 99801 162 99804
rect 810 99804 1584 99810
rect 810 99801 816 99804
rect 894 99764 900 99767
rect 126 99758 900 99764
rect 1548 99764 1554 99767
rect 1548 99758 1584 99764
rect 126 99724 138 99758
rect 1572 99724 1584 99758
rect 126 99718 900 99724
rect 894 99715 900 99718
rect 1548 99718 1584 99724
rect 1548 99715 1554 99718
rect 156 99678 162 99681
rect 126 99672 162 99678
rect 810 99678 816 99681
rect 810 99672 1584 99678
rect 126 99638 138 99672
rect 1572 99638 1584 99672
rect 126 99632 162 99638
rect 156 99629 162 99632
rect 810 99632 1584 99638
rect 810 99629 816 99632
rect 894 99592 900 99595
rect 126 99586 900 99592
rect 1548 99592 1554 99595
rect 1548 99586 1584 99592
rect 126 99552 138 99586
rect 1572 99552 1584 99586
rect 126 99546 900 99552
rect 894 99543 900 99546
rect 1548 99546 1584 99552
rect 1548 99543 1554 99546
rect 156 99506 162 99509
rect 126 99500 162 99506
rect 810 99506 816 99509
rect 810 99500 1584 99506
rect 126 99466 138 99500
rect 1572 99466 1584 99500
rect 126 99460 162 99466
rect 156 99457 162 99460
rect 810 99460 1584 99466
rect 810 99457 816 99460
rect 894 99420 900 99423
rect 126 99414 900 99420
rect 1548 99420 1554 99423
rect 1548 99414 1584 99420
rect 126 99380 138 99414
rect 1572 99380 1584 99414
rect 126 99374 900 99380
rect 894 99371 900 99374
rect 1548 99374 1584 99380
rect 1548 99371 1554 99374
rect 156 99334 162 99337
rect 126 99328 162 99334
rect 810 99334 816 99337
rect 810 99328 1584 99334
rect 126 99294 138 99328
rect 1572 99294 1584 99328
rect 126 99288 162 99294
rect 156 99285 162 99288
rect 810 99288 1584 99294
rect 810 99285 816 99288
rect 894 99248 900 99251
rect 126 99242 900 99248
rect 1548 99248 1554 99251
rect 1548 99242 1584 99248
rect 126 99208 138 99242
rect 1572 99208 1584 99242
rect 126 99202 900 99208
rect 894 99199 900 99202
rect 1548 99202 1584 99208
rect 1548 99199 1554 99202
rect 156 99162 162 99165
rect 126 99156 162 99162
rect 810 99162 816 99165
rect 810 99156 1584 99162
rect 126 99122 138 99156
rect 1572 99122 1584 99156
rect 126 99116 162 99122
rect 156 99113 162 99116
rect 810 99116 1584 99122
rect 810 99113 816 99116
rect 894 99076 900 99079
rect 126 99070 900 99076
rect 1548 99076 1554 99079
rect 1548 99070 1584 99076
rect 126 99036 138 99070
rect 1572 99036 1584 99070
rect 126 99030 900 99036
rect 894 99027 900 99030
rect 1548 99030 1584 99036
rect 1548 99027 1554 99030
rect 156 98990 162 98993
rect 126 98984 162 98990
rect 810 98990 816 98993
rect 810 98984 1584 98990
rect 126 98950 138 98984
rect 1572 98950 1584 98984
rect 126 98944 162 98950
rect 156 98941 162 98944
rect 810 98944 1584 98950
rect 810 98941 816 98944
rect 894 98904 900 98907
rect 126 98898 900 98904
rect 1548 98904 1554 98907
rect 1548 98898 1584 98904
rect 126 98864 138 98898
rect 1572 98864 1584 98898
rect 126 98858 900 98864
rect 894 98855 900 98858
rect 1548 98858 1584 98864
rect 1548 98855 1554 98858
rect 156 98818 162 98821
rect 126 98812 162 98818
rect 810 98818 816 98821
rect 810 98812 1584 98818
rect 126 98778 138 98812
rect 1572 98778 1584 98812
rect 126 98772 162 98778
rect 156 98769 162 98772
rect 810 98772 1584 98778
rect 810 98769 816 98772
rect 894 98732 900 98735
rect 126 98726 900 98732
rect 1548 98732 1554 98735
rect 1548 98726 1584 98732
rect 126 98692 138 98726
rect 1572 98692 1584 98726
rect 126 98686 900 98692
rect 894 98683 900 98686
rect 1548 98686 1584 98692
rect 1548 98683 1554 98686
rect 156 98646 162 98649
rect 126 98640 162 98646
rect 810 98646 816 98649
rect 810 98640 1584 98646
rect 126 98606 138 98640
rect 1572 98606 1584 98640
rect 126 98600 162 98606
rect 156 98597 162 98600
rect 810 98600 1584 98606
rect 810 98597 816 98600
rect 894 98560 900 98563
rect 126 98554 900 98560
rect 1548 98560 1554 98563
rect 1548 98554 1584 98560
rect 126 98520 138 98554
rect 1572 98520 1584 98554
rect 126 98514 900 98520
rect 894 98511 900 98514
rect 1548 98514 1584 98520
rect 1548 98511 1554 98514
rect 156 98474 162 98477
rect 126 98468 162 98474
rect 810 98474 816 98477
rect 810 98468 1584 98474
rect 126 98434 138 98468
rect 1572 98434 1584 98468
rect 126 98428 162 98434
rect 156 98425 162 98428
rect 810 98428 1584 98434
rect 810 98425 816 98428
rect 894 98388 900 98391
rect 126 98382 900 98388
rect 1548 98388 1554 98391
rect 1548 98382 1584 98388
rect 126 98348 138 98382
rect 1572 98348 1584 98382
rect 126 98342 900 98348
rect 894 98339 900 98342
rect 1548 98342 1584 98348
rect 1548 98339 1554 98342
rect 156 98302 162 98305
rect 126 98296 162 98302
rect 810 98302 816 98305
rect 810 98296 1584 98302
rect 126 98262 138 98296
rect 1572 98262 1584 98296
rect 126 98256 162 98262
rect 156 98253 162 98256
rect 810 98256 1584 98262
rect 810 98253 816 98256
rect 894 98216 900 98219
rect 126 98210 900 98216
rect 1548 98216 1554 98219
rect 1548 98210 1584 98216
rect 126 98176 138 98210
rect 1572 98176 1584 98210
rect 126 98170 900 98176
rect 894 98167 900 98170
rect 1548 98170 1584 98176
rect 1548 98167 1554 98170
rect 156 98130 162 98133
rect 126 98124 162 98130
rect 810 98130 816 98133
rect 810 98124 1584 98130
rect 126 98090 138 98124
rect 1572 98090 1584 98124
rect 126 98084 162 98090
rect 156 98081 162 98084
rect 810 98084 1584 98090
rect 810 98081 816 98084
rect 894 98044 900 98047
rect 126 98038 900 98044
rect 1548 98044 1554 98047
rect 1548 98038 1584 98044
rect 126 98004 138 98038
rect 1572 98004 1584 98038
rect 126 97998 900 98004
rect 894 97995 900 97998
rect 1548 97998 1584 98004
rect 1548 97995 1554 97998
rect 156 97958 162 97961
rect 126 97952 162 97958
rect 810 97958 816 97961
rect 810 97952 1584 97958
rect 126 97918 138 97952
rect 1572 97918 1584 97952
rect 126 97912 162 97918
rect 156 97909 162 97912
rect 810 97912 1584 97918
rect 810 97909 816 97912
rect 894 97872 900 97875
rect 126 97866 900 97872
rect 1548 97872 1554 97875
rect 1548 97866 1584 97872
rect 126 97832 138 97866
rect 1572 97832 1584 97866
rect 126 97826 900 97832
rect 894 97823 900 97826
rect 1548 97826 1584 97832
rect 1548 97823 1554 97826
rect 156 97786 162 97789
rect 126 97780 162 97786
rect 810 97786 816 97789
rect 810 97780 1584 97786
rect 126 97746 138 97780
rect 1572 97746 1584 97780
rect 126 97740 162 97746
rect 156 97737 162 97740
rect 810 97740 1584 97746
rect 810 97737 816 97740
rect 894 97700 900 97703
rect 126 97694 900 97700
rect 1548 97700 1554 97703
rect 1548 97694 1584 97700
rect 126 97660 138 97694
rect 1572 97660 1584 97694
rect 126 97654 900 97660
rect 894 97651 900 97654
rect 1548 97654 1584 97660
rect 1548 97651 1554 97654
rect 156 97614 162 97617
rect 126 97608 162 97614
rect 810 97614 816 97617
rect 810 97608 1584 97614
rect 126 97574 138 97608
rect 1572 97574 1584 97608
rect 126 97568 162 97574
rect 156 97565 162 97568
rect 810 97568 1584 97574
rect 810 97565 816 97568
rect 894 97528 900 97531
rect 126 97522 900 97528
rect 1548 97528 1554 97531
rect 1548 97522 1584 97528
rect 126 97488 138 97522
rect 1572 97488 1584 97522
rect 126 97482 900 97488
rect 894 97479 900 97482
rect 1548 97482 1584 97488
rect 1548 97479 1554 97482
rect 156 97442 162 97445
rect 126 97436 162 97442
rect 810 97442 816 97445
rect 810 97436 1584 97442
rect 126 97402 138 97436
rect 1572 97402 1584 97436
rect 126 97396 162 97402
rect 156 97393 162 97396
rect 810 97396 1584 97402
rect 810 97393 816 97396
rect 894 97356 900 97359
rect 126 97350 900 97356
rect 1548 97356 1554 97359
rect 1548 97350 1584 97356
rect 126 97316 138 97350
rect 1572 97316 1584 97350
rect 126 97310 900 97316
rect 894 97307 900 97310
rect 1548 97310 1584 97316
rect 1548 97307 1554 97310
rect 156 97270 162 97273
rect 126 97264 162 97270
rect 810 97270 816 97273
rect 810 97264 1584 97270
rect 126 97230 138 97264
rect 1572 97230 1584 97264
rect 126 97224 162 97230
rect 156 97221 162 97224
rect 810 97224 1584 97230
rect 810 97221 816 97224
rect 894 97184 900 97187
rect 126 97178 900 97184
rect 1548 97184 1554 97187
rect 1548 97178 1584 97184
rect 126 97144 138 97178
rect 1572 97144 1584 97178
rect 126 97138 900 97144
rect 894 97135 900 97138
rect 1548 97138 1584 97144
rect 1548 97135 1554 97138
rect 156 97098 162 97101
rect 126 97092 162 97098
rect 810 97098 816 97101
rect 810 97092 1584 97098
rect 126 97058 138 97092
rect 1572 97058 1584 97092
rect 126 97052 162 97058
rect 156 97049 162 97052
rect 810 97052 1584 97058
rect 810 97049 816 97052
rect 894 97012 900 97015
rect 126 97006 900 97012
rect 1548 97012 1554 97015
rect 1548 97006 1584 97012
rect 126 96972 138 97006
rect 1572 96972 1584 97006
rect 126 96966 900 96972
rect 894 96963 900 96966
rect 1548 96966 1584 96972
rect 1548 96963 1554 96966
rect 156 96926 162 96929
rect 126 96920 162 96926
rect 810 96926 816 96929
rect 810 96920 1584 96926
rect 126 96886 138 96920
rect 1572 96886 1584 96920
rect 126 96880 162 96886
rect 156 96877 162 96880
rect 810 96880 1584 96886
rect 810 96877 816 96880
rect 894 96840 900 96843
rect 126 96834 900 96840
rect 1548 96840 1554 96843
rect 1548 96834 1584 96840
rect 126 96800 138 96834
rect 1572 96800 1584 96834
rect 126 96794 900 96800
rect 894 96791 900 96794
rect 1548 96794 1584 96800
rect 1548 96791 1554 96794
rect 156 96754 162 96757
rect 126 96748 162 96754
rect 810 96754 816 96757
rect 810 96748 1584 96754
rect 126 96714 138 96748
rect 1572 96714 1584 96748
rect 126 96708 162 96714
rect 156 96705 162 96708
rect 810 96708 1584 96714
rect 810 96705 816 96708
rect 894 96668 900 96671
rect 126 96662 900 96668
rect 1548 96668 1554 96671
rect 1548 96662 1584 96668
rect 126 96628 138 96662
rect 1572 96628 1584 96662
rect 126 96622 900 96628
rect 894 96619 900 96622
rect 1548 96622 1584 96628
rect 1548 96619 1554 96622
rect 156 96582 162 96585
rect 126 96576 162 96582
rect 810 96582 816 96585
rect 810 96576 1584 96582
rect 126 96542 138 96576
rect 1572 96542 1584 96576
rect 126 96536 162 96542
rect 156 96533 162 96536
rect 810 96536 1584 96542
rect 810 96533 816 96536
rect 894 96496 900 96499
rect 126 96490 900 96496
rect 1548 96496 1554 96499
rect 1548 96490 1584 96496
rect 126 96456 138 96490
rect 1572 96456 1584 96490
rect 126 96450 900 96456
rect 894 96447 900 96450
rect 1548 96450 1584 96456
rect 1548 96447 1554 96450
rect 156 96410 162 96413
rect 126 96404 162 96410
rect 810 96410 816 96413
rect 810 96404 1584 96410
rect 126 96370 138 96404
rect 1572 96370 1584 96404
rect 126 96364 162 96370
rect 156 96361 162 96364
rect 810 96364 1584 96370
rect 810 96361 816 96364
rect 894 96324 900 96327
rect 126 96318 900 96324
rect 1548 96324 1554 96327
rect 1548 96318 1584 96324
rect 126 96284 138 96318
rect 1572 96284 1584 96318
rect 126 96278 900 96284
rect 894 96275 900 96278
rect 1548 96278 1584 96284
rect 1548 96275 1554 96278
rect 156 96238 162 96241
rect 126 96232 162 96238
rect 810 96238 816 96241
rect 810 96232 1584 96238
rect 126 96198 138 96232
rect 1572 96198 1584 96232
rect 126 96192 162 96198
rect 156 96189 162 96192
rect 810 96192 1584 96198
rect 810 96189 816 96192
rect 894 96152 900 96155
rect 126 96146 900 96152
rect 1548 96152 1554 96155
rect 1548 96146 1584 96152
rect 126 96112 138 96146
rect 1572 96112 1584 96146
rect 126 96106 900 96112
rect 894 96103 900 96106
rect 1548 96106 1584 96112
rect 1548 96103 1554 96106
rect 156 96066 162 96069
rect 126 96060 162 96066
rect 810 96066 816 96069
rect 810 96060 1584 96066
rect 126 96026 138 96060
rect 1572 96026 1584 96060
rect 126 96020 162 96026
rect 156 96017 162 96020
rect 810 96020 1584 96026
rect 810 96017 816 96020
rect 894 95980 900 95983
rect 126 95974 900 95980
rect 1548 95980 1554 95983
rect 1548 95974 1584 95980
rect 126 95940 138 95974
rect 1572 95940 1584 95974
rect 126 95934 900 95940
rect 894 95931 900 95934
rect 1548 95934 1584 95940
rect 1548 95931 1554 95934
rect 156 95894 162 95897
rect 126 95888 162 95894
rect 810 95894 816 95897
rect 810 95888 1584 95894
rect 126 95854 138 95888
rect 1572 95854 1584 95888
rect 126 95848 162 95854
rect 156 95845 162 95848
rect 810 95848 1584 95854
rect 810 95845 816 95848
rect 894 95808 900 95811
rect 126 95802 900 95808
rect 1548 95808 1554 95811
rect 1548 95802 1584 95808
rect 126 95768 138 95802
rect 1572 95768 1584 95802
rect 126 95762 900 95768
rect 894 95759 900 95762
rect 1548 95762 1584 95768
rect 1548 95759 1554 95762
rect 156 95722 162 95725
rect 126 95716 162 95722
rect 810 95722 816 95725
rect 810 95716 1584 95722
rect 126 95682 138 95716
rect 1572 95682 1584 95716
rect 126 95676 162 95682
rect 156 95673 162 95676
rect 810 95676 1584 95682
rect 810 95673 816 95676
rect 894 95636 900 95639
rect 126 95630 900 95636
rect 1548 95636 1554 95639
rect 1548 95630 1584 95636
rect 126 95596 138 95630
rect 1572 95596 1584 95630
rect 126 95590 900 95596
rect 894 95587 900 95590
rect 1548 95590 1584 95596
rect 1548 95587 1554 95590
rect 156 95550 162 95553
rect 126 95544 162 95550
rect 810 95550 816 95553
rect 810 95544 1584 95550
rect 126 95510 138 95544
rect 1572 95510 1584 95544
rect 126 95504 162 95510
rect 156 95501 162 95504
rect 810 95504 1584 95510
rect 810 95501 816 95504
rect 894 95464 900 95467
rect 126 95458 900 95464
rect 1548 95464 1554 95467
rect 1548 95458 1584 95464
rect 126 95424 138 95458
rect 1572 95424 1584 95458
rect 126 95418 900 95424
rect 894 95415 900 95418
rect 1548 95418 1584 95424
rect 1548 95415 1554 95418
rect 156 95378 162 95381
rect 126 95372 162 95378
rect 810 95378 816 95381
rect 810 95372 1584 95378
rect 126 95338 138 95372
rect 1572 95338 1584 95372
rect 126 95332 162 95338
rect 156 95329 162 95332
rect 810 95332 1584 95338
rect 810 95329 816 95332
rect 894 95292 900 95295
rect 126 95286 900 95292
rect 1548 95292 1554 95295
rect 1548 95286 1584 95292
rect 126 95252 138 95286
rect 1572 95252 1584 95286
rect 126 95246 900 95252
rect 894 95243 900 95246
rect 1548 95246 1584 95252
rect 1548 95243 1554 95246
rect 156 95206 162 95209
rect 126 95200 162 95206
rect 810 95206 816 95209
rect 810 95200 1584 95206
rect 126 95166 138 95200
rect 1572 95166 1584 95200
rect 126 95160 162 95166
rect 156 95157 162 95160
rect 810 95160 1584 95166
rect 810 95157 816 95160
rect 894 95120 900 95123
rect 126 95114 900 95120
rect 1548 95120 1554 95123
rect 1548 95114 1584 95120
rect 126 95080 138 95114
rect 1572 95080 1584 95114
rect 126 95074 900 95080
rect 894 95071 900 95074
rect 1548 95074 1584 95080
rect 1548 95071 1554 95074
rect 156 95034 162 95037
rect 126 95028 162 95034
rect 810 95034 816 95037
rect 810 95028 1584 95034
rect 126 94994 138 95028
rect 1572 94994 1584 95028
rect 126 94988 162 94994
rect 156 94985 162 94988
rect 810 94988 1584 94994
rect 810 94985 816 94988
rect 894 94948 900 94951
rect 126 94942 900 94948
rect 1548 94948 1554 94951
rect 1548 94942 1584 94948
rect 126 94908 138 94942
rect 1572 94908 1584 94942
rect 126 94902 900 94908
rect 894 94899 900 94902
rect 1548 94902 1584 94908
rect 1548 94899 1554 94902
rect 156 94862 162 94865
rect 126 94856 162 94862
rect 810 94862 816 94865
rect 810 94856 1584 94862
rect 126 94822 138 94856
rect 1572 94822 1584 94856
rect 126 94816 162 94822
rect 156 94813 162 94816
rect 810 94816 1584 94822
rect 810 94813 816 94816
rect 894 94776 900 94779
rect 126 94770 900 94776
rect 1548 94776 1554 94779
rect 1548 94770 1584 94776
rect 126 94736 138 94770
rect 1572 94736 1584 94770
rect 126 94730 900 94736
rect 894 94727 900 94730
rect 1548 94730 1584 94736
rect 1548 94727 1554 94730
rect 156 94690 162 94693
rect 126 94684 162 94690
rect 810 94690 816 94693
rect 810 94684 1584 94690
rect 126 94650 138 94684
rect 1572 94650 1584 94684
rect 126 94644 162 94650
rect 156 94641 162 94644
rect 810 94644 1584 94650
rect 810 94641 816 94644
rect 894 94604 900 94607
rect 126 94598 900 94604
rect 1548 94604 1554 94607
rect 1548 94598 1584 94604
rect 126 94564 138 94598
rect 1572 94564 1584 94598
rect 126 94558 900 94564
rect 894 94555 900 94558
rect 1548 94558 1584 94564
rect 1548 94555 1554 94558
rect 156 94518 162 94521
rect 126 94512 162 94518
rect 810 94518 816 94521
rect 810 94512 1584 94518
rect 126 94478 138 94512
rect 1572 94478 1584 94512
rect 126 94472 162 94478
rect 156 94469 162 94472
rect 810 94472 1584 94478
rect 810 94469 816 94472
rect 894 94432 900 94435
rect 126 94426 900 94432
rect 1548 94432 1554 94435
rect 1548 94426 1584 94432
rect 126 94392 138 94426
rect 1572 94392 1584 94426
rect 126 94386 900 94392
rect 894 94383 900 94386
rect 1548 94386 1584 94392
rect 1548 94383 1554 94386
rect 156 94346 162 94349
rect 126 94340 162 94346
rect 810 94346 816 94349
rect 810 94340 1584 94346
rect 126 94306 138 94340
rect 1572 94306 1584 94340
rect 126 94300 162 94306
rect 156 94297 162 94300
rect 810 94300 1584 94306
rect 810 94297 816 94300
rect 894 94260 900 94263
rect 126 94254 900 94260
rect 1548 94260 1554 94263
rect 1548 94254 1584 94260
rect 126 94220 138 94254
rect 1572 94220 1584 94254
rect 126 94214 900 94220
rect 894 94211 900 94214
rect 1548 94214 1584 94220
rect 1548 94211 1554 94214
rect 156 94174 162 94177
rect 126 94168 162 94174
rect 810 94174 816 94177
rect 810 94168 1584 94174
rect 126 94134 138 94168
rect 1572 94134 1584 94168
rect 126 94128 162 94134
rect 156 94125 162 94128
rect 810 94128 1584 94134
rect 810 94125 816 94128
rect 894 94088 900 94091
rect 126 94082 900 94088
rect 1548 94088 1554 94091
rect 1548 94082 1584 94088
rect 126 94048 138 94082
rect 1572 94048 1584 94082
rect 126 94042 900 94048
rect 894 94039 900 94042
rect 1548 94042 1584 94048
rect 1548 94039 1554 94042
rect 156 94002 162 94005
rect 126 93996 162 94002
rect 810 94002 816 94005
rect 810 93996 1584 94002
rect 126 93962 138 93996
rect 1572 93962 1584 93996
rect 126 93956 162 93962
rect 156 93953 162 93956
rect 810 93956 1584 93962
rect 810 93953 816 93956
rect 894 93916 900 93919
rect 126 93910 900 93916
rect 1548 93916 1554 93919
rect 1548 93910 1584 93916
rect 126 93876 138 93910
rect 1572 93876 1584 93910
rect 126 93870 900 93876
rect 894 93867 900 93870
rect 1548 93870 1584 93876
rect 1548 93867 1554 93870
rect 156 93830 162 93833
rect 126 93824 162 93830
rect 810 93830 816 93833
rect 810 93824 1584 93830
rect 126 93790 138 93824
rect 1572 93790 1584 93824
rect 126 93784 162 93790
rect 156 93781 162 93784
rect 810 93784 1584 93790
rect 810 93781 816 93784
rect 894 93744 900 93747
rect 126 93738 900 93744
rect 1548 93744 1554 93747
rect 1548 93738 1584 93744
rect 126 93704 138 93738
rect 1572 93704 1584 93738
rect 126 93698 900 93704
rect 894 93695 900 93698
rect 1548 93698 1584 93704
rect 1548 93695 1554 93698
rect 156 93658 162 93661
rect 126 93652 162 93658
rect 810 93658 816 93661
rect 810 93652 1584 93658
rect 126 93618 138 93652
rect 1572 93618 1584 93652
rect 126 93612 162 93618
rect 156 93609 162 93612
rect 810 93612 1584 93618
rect 810 93609 816 93612
rect 894 93572 900 93575
rect 126 93566 900 93572
rect 1548 93572 1554 93575
rect 1548 93566 1584 93572
rect 126 93532 138 93566
rect 1572 93532 1584 93566
rect 126 93526 900 93532
rect 894 93523 900 93526
rect 1548 93526 1584 93532
rect 1548 93523 1554 93526
rect 156 93486 162 93489
rect 126 93480 162 93486
rect 810 93486 816 93489
rect 810 93480 1584 93486
rect 126 93446 138 93480
rect 1572 93446 1584 93480
rect 126 93440 162 93446
rect 156 93437 162 93440
rect 810 93440 1584 93446
rect 810 93437 816 93440
rect 894 93400 900 93403
rect 126 93394 900 93400
rect 1548 93400 1554 93403
rect 1548 93394 1584 93400
rect 126 93360 138 93394
rect 1572 93360 1584 93394
rect 126 93354 900 93360
rect 894 93351 900 93354
rect 1548 93354 1584 93360
rect 1548 93351 1554 93354
rect 156 93314 162 93317
rect 126 93308 162 93314
rect 810 93314 816 93317
rect 810 93308 1584 93314
rect 126 93274 138 93308
rect 1572 93274 1584 93308
rect 126 93268 162 93274
rect 156 93265 162 93268
rect 810 93268 1584 93274
rect 810 93265 816 93268
rect 894 93228 900 93231
rect 126 93222 900 93228
rect 1548 93228 1554 93231
rect 1548 93222 1584 93228
rect 126 93188 138 93222
rect 1572 93188 1584 93222
rect 126 93182 900 93188
rect 894 93179 900 93182
rect 1548 93182 1584 93188
rect 1548 93179 1554 93182
rect 156 93142 162 93145
rect 126 93136 162 93142
rect 810 93142 816 93145
rect 810 93136 1584 93142
rect 126 93102 138 93136
rect 1572 93102 1584 93136
rect 126 93096 162 93102
rect 156 93093 162 93096
rect 810 93096 1584 93102
rect 810 93093 816 93096
rect 894 93056 900 93059
rect 126 93050 900 93056
rect 1548 93056 1554 93059
rect 1548 93050 1584 93056
rect 126 93016 138 93050
rect 1572 93016 1584 93050
rect 126 93010 900 93016
rect 894 93007 900 93010
rect 1548 93010 1584 93016
rect 1548 93007 1554 93010
rect 156 92970 162 92973
rect 126 92964 162 92970
rect 810 92970 816 92973
rect 810 92964 1584 92970
rect 126 92930 138 92964
rect 1572 92930 1584 92964
rect 126 92924 162 92930
rect 156 92921 162 92924
rect 810 92924 1584 92930
rect 810 92921 816 92924
rect 894 92884 900 92887
rect 126 92878 900 92884
rect 1548 92884 1554 92887
rect 1548 92878 1584 92884
rect 126 92844 138 92878
rect 1572 92844 1584 92878
rect 126 92838 900 92844
rect 894 92835 900 92838
rect 1548 92838 1584 92844
rect 1548 92835 1554 92838
rect 156 92798 162 92801
rect 126 92792 162 92798
rect 810 92798 816 92801
rect 810 92792 1584 92798
rect 126 92758 138 92792
rect 1572 92758 1584 92792
rect 126 92752 162 92758
rect 156 92749 162 92752
rect 810 92752 1584 92758
rect 810 92749 816 92752
rect 894 92712 900 92715
rect 126 92706 900 92712
rect 1548 92712 1554 92715
rect 1548 92706 1584 92712
rect 126 92672 138 92706
rect 1572 92672 1584 92706
rect 126 92666 900 92672
rect 894 92663 900 92666
rect 1548 92666 1584 92672
rect 1548 92663 1554 92666
rect 156 92626 162 92629
rect 126 92620 162 92626
rect 810 92626 816 92629
rect 810 92620 1584 92626
rect 126 92586 138 92620
rect 1572 92586 1584 92620
rect 126 92580 162 92586
rect 156 92577 162 92580
rect 810 92580 1584 92586
rect 810 92577 816 92580
rect 894 92540 900 92543
rect 126 92534 900 92540
rect 1548 92540 1554 92543
rect 1548 92534 1584 92540
rect 126 92500 138 92534
rect 1572 92500 1584 92534
rect 126 92494 900 92500
rect 894 92491 900 92494
rect 1548 92494 1584 92500
rect 1548 92491 1554 92494
rect 156 92454 162 92457
rect 126 92448 162 92454
rect 810 92454 816 92457
rect 810 92448 1584 92454
rect 126 92414 138 92448
rect 1572 92414 1584 92448
rect 126 92408 162 92414
rect 156 92405 162 92408
rect 810 92408 1584 92414
rect 810 92405 816 92408
rect 894 92368 900 92371
rect 126 92362 900 92368
rect 1548 92368 1554 92371
rect 1548 92362 1584 92368
rect 126 92328 138 92362
rect 1572 92328 1584 92362
rect 126 92322 900 92328
rect 894 92319 900 92322
rect 1548 92322 1584 92328
rect 1548 92319 1554 92322
rect 156 92282 162 92285
rect 126 92276 162 92282
rect 810 92282 816 92285
rect 810 92276 1584 92282
rect 126 92242 138 92276
rect 1572 92242 1584 92276
rect 126 92236 162 92242
rect 156 92233 162 92236
rect 810 92236 1584 92242
rect 810 92233 816 92236
rect 894 92196 900 92199
rect 126 92190 900 92196
rect 1548 92196 1554 92199
rect 1548 92190 1584 92196
rect 126 92156 138 92190
rect 1572 92156 1584 92190
rect 126 92150 900 92156
rect 894 92147 900 92150
rect 1548 92150 1584 92156
rect 1548 92147 1554 92150
rect 156 92110 162 92113
rect 126 92104 162 92110
rect 810 92110 816 92113
rect 810 92104 1584 92110
rect 126 92070 138 92104
rect 1572 92070 1584 92104
rect 126 92064 162 92070
rect 156 92061 162 92064
rect 810 92064 1584 92070
rect 810 92061 816 92064
rect 894 92024 900 92027
rect 126 92018 900 92024
rect 1548 92024 1554 92027
rect 1548 92018 1584 92024
rect 126 91984 138 92018
rect 1572 91984 1584 92018
rect 126 91978 900 91984
rect 894 91975 900 91978
rect 1548 91978 1584 91984
rect 1548 91975 1554 91978
rect 156 91938 162 91941
rect 126 91932 162 91938
rect 810 91938 816 91941
rect 810 91932 1584 91938
rect 126 91898 138 91932
rect 1572 91898 1584 91932
rect 126 91892 162 91898
rect 156 91889 162 91892
rect 810 91892 1584 91898
rect 810 91889 816 91892
rect 894 91852 900 91855
rect 126 91846 900 91852
rect 1548 91852 1554 91855
rect 1548 91846 1584 91852
rect 126 91812 138 91846
rect 1572 91812 1584 91846
rect 126 91806 900 91812
rect 894 91803 900 91806
rect 1548 91806 1584 91812
rect 1548 91803 1554 91806
rect 156 91766 162 91769
rect 126 91760 162 91766
rect 810 91766 816 91769
rect 810 91760 1584 91766
rect 126 91726 138 91760
rect 1572 91726 1584 91760
rect 126 91720 162 91726
rect 156 91717 162 91720
rect 810 91720 1584 91726
rect 810 91717 816 91720
rect 894 91680 900 91683
rect 126 91674 900 91680
rect 1548 91680 1554 91683
rect 1548 91674 1584 91680
rect 126 91640 138 91674
rect 1572 91640 1584 91674
rect 126 91634 900 91640
rect 894 91631 900 91634
rect 1548 91634 1584 91640
rect 1548 91631 1554 91634
rect 156 91594 162 91597
rect 126 91588 162 91594
rect 810 91594 816 91597
rect 810 91588 1584 91594
rect 126 91554 138 91588
rect 1572 91554 1584 91588
rect 126 91548 162 91554
rect 156 91545 162 91548
rect 810 91548 1584 91554
rect 810 91545 816 91548
rect 894 91508 900 91511
rect 126 91502 900 91508
rect 1548 91508 1554 91511
rect 1548 91502 1584 91508
rect 126 91468 138 91502
rect 1572 91468 1584 91502
rect 126 91462 900 91468
rect 894 91459 900 91462
rect 1548 91462 1584 91468
rect 1548 91459 1554 91462
rect 156 91422 162 91425
rect 126 91416 162 91422
rect 810 91422 816 91425
rect 810 91416 1584 91422
rect 126 91382 138 91416
rect 1572 91382 1584 91416
rect 126 91376 162 91382
rect 156 91373 162 91376
rect 810 91376 1584 91382
rect 810 91373 816 91376
rect 894 91336 900 91339
rect 126 91330 900 91336
rect 1548 91336 1554 91339
rect 1548 91330 1584 91336
rect 126 91296 138 91330
rect 1572 91296 1584 91330
rect 126 91290 900 91296
rect 894 91287 900 91290
rect 1548 91290 1584 91296
rect 1548 91287 1554 91290
rect 156 91250 162 91253
rect 126 91244 162 91250
rect 810 91250 816 91253
rect 810 91244 1584 91250
rect 126 91210 138 91244
rect 1572 91210 1584 91244
rect 126 91204 162 91210
rect 156 91201 162 91204
rect 810 91204 1584 91210
rect 810 91201 816 91204
rect 894 91164 900 91167
rect 126 91158 900 91164
rect 1548 91164 1554 91167
rect 1548 91158 1584 91164
rect 126 91124 138 91158
rect 1572 91124 1584 91158
rect 126 91118 900 91124
rect 894 91115 900 91118
rect 1548 91118 1584 91124
rect 1548 91115 1554 91118
rect 156 91078 162 91081
rect 126 91072 162 91078
rect 810 91078 816 91081
rect 810 91072 1584 91078
rect 126 91038 138 91072
rect 1572 91038 1584 91072
rect 126 91032 162 91038
rect 156 91029 162 91032
rect 810 91032 1584 91038
rect 810 91029 816 91032
rect 894 90992 900 90995
rect 126 90986 900 90992
rect 1548 90992 1554 90995
rect 1548 90986 1584 90992
rect 126 90952 138 90986
rect 1572 90952 1584 90986
rect 126 90946 900 90952
rect 894 90943 900 90946
rect 1548 90946 1584 90952
rect 1548 90943 1554 90946
rect 156 90906 162 90909
rect 126 90900 162 90906
rect 810 90906 816 90909
rect 810 90900 1584 90906
rect 126 90866 138 90900
rect 1572 90866 1584 90900
rect 126 90860 162 90866
rect 156 90857 162 90860
rect 810 90860 1584 90866
rect 810 90857 816 90860
rect 894 90820 900 90823
rect 126 90814 900 90820
rect 1548 90820 1554 90823
rect 1548 90814 1584 90820
rect 126 90780 138 90814
rect 1572 90780 1584 90814
rect 126 90774 900 90780
rect 894 90771 900 90774
rect 1548 90774 1584 90780
rect 1548 90771 1554 90774
rect 156 90734 162 90737
rect 126 90728 162 90734
rect 810 90734 816 90737
rect 810 90728 1584 90734
rect 126 90694 138 90728
rect 1572 90694 1584 90728
rect 126 90688 162 90694
rect 156 90685 162 90688
rect 810 90688 1584 90694
rect 810 90685 816 90688
rect 894 90648 900 90651
rect 126 90642 900 90648
rect 1548 90648 1554 90651
rect 1548 90642 1584 90648
rect 126 90608 138 90642
rect 1572 90608 1584 90642
rect 126 90602 900 90608
rect 894 90599 900 90602
rect 1548 90602 1584 90608
rect 1548 90599 1554 90602
rect 156 90562 162 90565
rect 126 90556 162 90562
rect 810 90562 816 90565
rect 810 90556 1584 90562
rect 126 90522 138 90556
rect 1572 90522 1584 90556
rect 126 90516 162 90522
rect 156 90513 162 90516
rect 810 90516 1584 90522
rect 810 90513 816 90516
rect 894 90476 900 90479
rect 126 90470 900 90476
rect 1548 90476 1554 90479
rect 1548 90470 1584 90476
rect 126 90436 138 90470
rect 1572 90436 1584 90470
rect 126 90430 900 90436
rect 894 90427 900 90430
rect 1548 90430 1584 90436
rect 1548 90427 1554 90430
rect 156 90390 162 90393
rect 126 90384 162 90390
rect 810 90390 816 90393
rect 810 90384 1584 90390
rect 126 90350 138 90384
rect 1572 90350 1584 90384
rect 126 90344 162 90350
rect 156 90341 162 90344
rect 810 90344 1584 90350
rect 810 90341 816 90344
rect 894 90304 900 90307
rect 126 90298 900 90304
rect 1548 90304 1554 90307
rect 1548 90298 1584 90304
rect 126 90264 138 90298
rect 1572 90264 1584 90298
rect 126 90258 900 90264
rect 894 90255 900 90258
rect 1548 90258 1584 90264
rect 1548 90255 1554 90258
rect 156 90218 162 90221
rect 126 90212 162 90218
rect 810 90218 816 90221
rect 810 90212 1584 90218
rect 126 90178 138 90212
rect 1572 90178 1584 90212
rect 126 90172 162 90178
rect 156 90169 162 90172
rect 810 90172 1584 90178
rect 810 90169 816 90172
rect 894 90132 900 90135
rect 126 90126 900 90132
rect 1548 90132 1554 90135
rect 1548 90126 1584 90132
rect 126 90092 138 90126
rect 1572 90092 1584 90126
rect 126 90086 900 90092
rect 894 90083 900 90086
rect 1548 90086 1584 90092
rect 1548 90083 1554 90086
rect 156 90046 162 90049
rect 126 90040 162 90046
rect 810 90046 816 90049
rect 810 90040 1584 90046
rect 126 90006 138 90040
rect 1572 90006 1584 90040
rect 126 90000 162 90006
rect 156 89997 162 90000
rect 810 90000 1584 90006
rect 810 89997 816 90000
rect 894 89960 900 89963
rect 126 89954 900 89960
rect 1548 89960 1554 89963
rect 1548 89954 1584 89960
rect 126 89920 138 89954
rect 1572 89920 1584 89954
rect 126 89914 900 89920
rect 894 89911 900 89914
rect 1548 89914 1584 89920
rect 1548 89911 1554 89914
rect 156 89874 162 89877
rect 126 89868 162 89874
rect 810 89874 816 89877
rect 810 89868 1584 89874
rect 126 89834 138 89868
rect 1572 89834 1584 89868
rect 126 89828 162 89834
rect 156 89825 162 89828
rect 810 89828 1584 89834
rect 810 89825 816 89828
rect 894 89788 900 89791
rect 126 89782 900 89788
rect 1548 89788 1554 89791
rect 1548 89782 1584 89788
rect 126 89748 138 89782
rect 1572 89748 1584 89782
rect 126 89742 900 89748
rect 894 89739 900 89742
rect 1548 89742 1584 89748
rect 1548 89739 1554 89742
rect 156 89702 162 89705
rect 126 89696 162 89702
rect 810 89702 816 89705
rect 810 89696 1584 89702
rect 126 89662 138 89696
rect 1572 89662 1584 89696
rect 126 89656 162 89662
rect 156 89653 162 89656
rect 810 89656 1584 89662
rect 810 89653 816 89656
rect 894 89616 900 89619
rect 126 89610 900 89616
rect 1548 89616 1554 89619
rect 1548 89610 1584 89616
rect 126 89576 138 89610
rect 1572 89576 1584 89610
rect 126 89570 900 89576
rect 894 89567 900 89570
rect 1548 89570 1584 89576
rect 1548 89567 1554 89570
rect 156 89530 162 89533
rect 126 89524 162 89530
rect 810 89530 816 89533
rect 810 89524 1584 89530
rect 126 89490 138 89524
rect 1572 89490 1584 89524
rect 126 89484 162 89490
rect 156 89481 162 89484
rect 810 89484 1584 89490
rect 810 89481 816 89484
rect 894 89444 900 89447
rect 126 89438 900 89444
rect 1548 89444 1554 89447
rect 1548 89438 1584 89444
rect 126 89404 138 89438
rect 1572 89404 1584 89438
rect 126 89398 900 89404
rect 894 89395 900 89398
rect 1548 89398 1584 89404
rect 1548 89395 1554 89398
rect 156 89358 162 89361
rect 126 89352 162 89358
rect 810 89358 816 89361
rect 810 89352 1584 89358
rect 126 89318 138 89352
rect 1572 89318 1584 89352
rect 126 89312 162 89318
rect 156 89309 162 89312
rect 810 89312 1584 89318
rect 810 89309 816 89312
rect 894 89272 900 89275
rect 126 89266 900 89272
rect 1548 89272 1554 89275
rect 1548 89266 1584 89272
rect 126 89232 138 89266
rect 1572 89232 1584 89266
rect 126 89226 900 89232
rect 894 89223 900 89226
rect 1548 89226 1584 89232
rect 1548 89223 1554 89226
rect 156 89186 162 89189
rect 126 89180 162 89186
rect 810 89186 816 89189
rect 810 89180 1584 89186
rect 126 89146 138 89180
rect 1572 89146 1584 89180
rect 126 89140 162 89146
rect 156 89137 162 89140
rect 810 89140 1584 89146
rect 810 89137 816 89140
rect 894 89100 900 89103
rect 126 89094 900 89100
rect 1548 89100 1554 89103
rect 1548 89094 1584 89100
rect 126 89060 138 89094
rect 1572 89060 1584 89094
rect 126 89054 900 89060
rect 894 89051 900 89054
rect 1548 89054 1584 89060
rect 1548 89051 1554 89054
rect 156 89014 162 89017
rect 126 89008 162 89014
rect 810 89014 816 89017
rect 810 89008 1584 89014
rect 126 88974 138 89008
rect 1572 88974 1584 89008
rect 126 88968 162 88974
rect 156 88965 162 88968
rect 810 88968 1584 88974
rect 810 88965 816 88968
rect 894 88928 900 88931
rect 126 88922 900 88928
rect 1548 88928 1554 88931
rect 1548 88922 1584 88928
rect 126 88888 138 88922
rect 1572 88888 1584 88922
rect 126 88882 900 88888
rect 894 88879 900 88882
rect 1548 88882 1584 88888
rect 1548 88879 1554 88882
rect 156 88842 162 88845
rect 126 88836 162 88842
rect 810 88842 816 88845
rect 810 88836 1584 88842
rect 126 88802 138 88836
rect 1572 88802 1584 88836
rect 126 88796 162 88802
rect 156 88793 162 88796
rect 810 88796 1584 88802
rect 810 88793 816 88796
rect 894 88756 900 88759
rect 126 88750 900 88756
rect 1548 88756 1554 88759
rect 1548 88750 1584 88756
rect 126 88716 138 88750
rect 1572 88716 1584 88750
rect 126 88710 900 88716
rect 894 88707 900 88710
rect 1548 88710 1584 88716
rect 1548 88707 1554 88710
rect 156 88670 162 88673
rect 126 88664 162 88670
rect 810 88670 816 88673
rect 810 88664 1584 88670
rect 126 88630 138 88664
rect 1572 88630 1584 88664
rect 126 88624 162 88630
rect 156 88621 162 88624
rect 810 88624 1584 88630
rect 810 88621 816 88624
rect 894 88584 900 88587
rect 126 88578 900 88584
rect 1548 88584 1554 88587
rect 1548 88578 1584 88584
rect 126 88544 138 88578
rect 1572 88544 1584 88578
rect 126 88538 900 88544
rect 894 88535 900 88538
rect 1548 88538 1584 88544
rect 1548 88535 1554 88538
rect 156 88498 162 88501
rect 126 88492 162 88498
rect 810 88498 816 88501
rect 810 88492 1584 88498
rect 126 88458 138 88492
rect 1572 88458 1584 88492
rect 126 88452 162 88458
rect 156 88449 162 88452
rect 810 88452 1584 88458
rect 810 88449 816 88452
rect 894 88412 900 88415
rect 126 88406 900 88412
rect 1548 88412 1554 88415
rect 1548 88406 1584 88412
rect 126 88372 138 88406
rect 1572 88372 1584 88406
rect 126 88366 900 88372
rect 894 88363 900 88366
rect 1548 88366 1584 88372
rect 1548 88363 1554 88366
rect 156 88326 162 88329
rect 126 88320 162 88326
rect 810 88326 816 88329
rect 810 88320 1584 88326
rect 126 88286 138 88320
rect 1572 88286 1584 88320
rect 126 88280 162 88286
rect 156 88277 162 88280
rect 810 88280 1584 88286
rect 810 88277 816 88280
rect 894 88240 900 88243
rect 126 88234 900 88240
rect 1548 88240 1554 88243
rect 1548 88234 1584 88240
rect 126 88200 138 88234
rect 1572 88200 1584 88234
rect 126 88194 900 88200
rect 894 88191 900 88194
rect 1548 88194 1584 88200
rect 1548 88191 1554 88194
rect 156 88154 162 88157
rect 126 88148 162 88154
rect 810 88154 816 88157
rect 810 88148 1584 88154
rect 126 88114 138 88148
rect 1572 88114 1584 88148
rect 126 88108 162 88114
rect 156 88105 162 88108
rect 810 88108 1584 88114
rect 810 88105 816 88108
rect 894 88068 900 88071
rect 126 88062 900 88068
rect 1548 88068 1554 88071
rect 1548 88062 1584 88068
rect 126 88028 138 88062
rect 1572 88028 1584 88062
rect 126 88022 900 88028
rect 894 88019 900 88022
rect 1548 88022 1584 88028
rect 1548 88019 1554 88022
rect 156 87982 162 87985
rect 126 87976 162 87982
rect 810 87982 816 87985
rect 810 87976 1584 87982
rect 126 87942 138 87976
rect 1572 87942 1584 87976
rect 126 87936 162 87942
rect 156 87933 162 87936
rect 810 87936 1584 87942
rect 810 87933 816 87936
rect 894 87896 900 87899
rect 126 87890 900 87896
rect 1548 87896 1554 87899
rect 1548 87890 1584 87896
rect 126 87856 138 87890
rect 1572 87856 1584 87890
rect 126 87850 900 87856
rect 894 87847 900 87850
rect 1548 87850 1584 87856
rect 1548 87847 1554 87850
rect 156 87810 162 87813
rect 126 87804 162 87810
rect 810 87810 816 87813
rect 810 87804 1584 87810
rect 126 87770 138 87804
rect 1572 87770 1584 87804
rect 126 87764 162 87770
rect 156 87761 162 87764
rect 810 87764 1584 87770
rect 810 87761 816 87764
rect 894 87724 900 87727
rect 126 87718 900 87724
rect 1548 87724 1554 87727
rect 1548 87718 1584 87724
rect 126 87684 138 87718
rect 1572 87684 1584 87718
rect 126 87678 900 87684
rect 894 87675 900 87678
rect 1548 87678 1584 87684
rect 1548 87675 1554 87678
rect 156 87638 162 87641
rect 126 87632 162 87638
rect 810 87638 816 87641
rect 810 87632 1584 87638
rect 126 87598 138 87632
rect 1572 87598 1584 87632
rect 126 87592 162 87598
rect 156 87589 162 87592
rect 810 87592 1584 87598
rect 810 87589 816 87592
rect 894 87552 900 87555
rect 126 87546 900 87552
rect 1548 87552 1554 87555
rect 1548 87546 1584 87552
rect 126 87512 138 87546
rect 1572 87512 1584 87546
rect 126 87506 900 87512
rect 894 87503 900 87506
rect 1548 87506 1584 87512
rect 1548 87503 1554 87506
rect 156 87466 162 87469
rect 126 87460 162 87466
rect 810 87466 816 87469
rect 810 87460 1584 87466
rect 126 87426 138 87460
rect 1572 87426 1584 87460
rect 126 87420 162 87426
rect 156 87417 162 87420
rect 810 87420 1584 87426
rect 810 87417 816 87420
rect 894 87380 900 87383
rect 126 87374 900 87380
rect 1548 87380 1554 87383
rect 1548 87374 1584 87380
rect 126 87340 138 87374
rect 1572 87340 1584 87374
rect 126 87334 900 87340
rect 894 87331 900 87334
rect 1548 87334 1584 87340
rect 1548 87331 1554 87334
rect 156 87294 162 87297
rect 126 87288 162 87294
rect 810 87294 816 87297
rect 810 87288 1584 87294
rect 126 87254 138 87288
rect 1572 87254 1584 87288
rect 126 87248 162 87254
rect 156 87245 162 87248
rect 810 87248 1584 87254
rect 810 87245 816 87248
rect 894 87208 900 87211
rect 126 87202 900 87208
rect 1548 87208 1554 87211
rect 1548 87202 1584 87208
rect 126 87168 138 87202
rect 1572 87168 1584 87202
rect 126 87162 900 87168
rect 894 87159 900 87162
rect 1548 87162 1584 87168
rect 1548 87159 1554 87162
rect 156 87122 162 87125
rect 126 87116 162 87122
rect 810 87122 816 87125
rect 810 87116 1584 87122
rect 126 87082 138 87116
rect 1572 87082 1584 87116
rect 126 87076 162 87082
rect 156 87073 162 87076
rect 810 87076 1584 87082
rect 810 87073 816 87076
rect 894 87036 900 87039
rect 126 87030 900 87036
rect 1548 87036 1554 87039
rect 1548 87030 1584 87036
rect 126 86996 138 87030
rect 1572 86996 1584 87030
rect 126 86990 900 86996
rect 894 86987 900 86990
rect 1548 86990 1584 86996
rect 1548 86987 1554 86990
rect 156 86950 162 86953
rect 126 86944 162 86950
rect 810 86950 816 86953
rect 810 86944 1584 86950
rect 126 86910 138 86944
rect 1572 86910 1584 86944
rect 126 86904 162 86910
rect 156 86901 162 86904
rect 810 86904 1584 86910
rect 810 86901 816 86904
rect 894 86864 900 86867
rect 126 86858 900 86864
rect 1548 86864 1554 86867
rect 1548 86858 1584 86864
rect 126 86824 138 86858
rect 1572 86824 1584 86858
rect 126 86818 900 86824
rect 894 86815 900 86818
rect 1548 86818 1584 86824
rect 1548 86815 1554 86818
rect 156 86778 162 86781
rect 126 86772 162 86778
rect 810 86778 816 86781
rect 810 86772 1584 86778
rect 126 86738 138 86772
rect 1572 86738 1584 86772
rect 126 86732 162 86738
rect 156 86729 162 86732
rect 810 86732 1584 86738
rect 810 86729 816 86732
rect 894 86692 900 86695
rect 126 86686 900 86692
rect 1548 86692 1554 86695
rect 1548 86686 1584 86692
rect 126 86652 138 86686
rect 1572 86652 1584 86686
rect 126 86646 900 86652
rect 894 86643 900 86646
rect 1548 86646 1584 86652
rect 1548 86643 1554 86646
rect 156 86606 162 86609
rect 126 86600 162 86606
rect 810 86606 816 86609
rect 810 86600 1584 86606
rect 126 86566 138 86600
rect 1572 86566 1584 86600
rect 126 86560 162 86566
rect 156 86557 162 86560
rect 810 86560 1584 86566
rect 810 86557 816 86560
rect 894 86520 900 86523
rect 126 86514 900 86520
rect 1548 86520 1554 86523
rect 1548 86514 1584 86520
rect 126 86480 138 86514
rect 1572 86480 1584 86514
rect 126 86474 900 86480
rect 894 86471 900 86474
rect 1548 86474 1584 86480
rect 1548 86471 1554 86474
rect 156 86434 162 86437
rect 126 86428 162 86434
rect 810 86434 816 86437
rect 810 86428 1584 86434
rect 126 86394 138 86428
rect 1572 86394 1584 86428
rect 126 86388 162 86394
rect 156 86385 162 86388
rect 810 86388 1584 86394
rect 810 86385 816 86388
rect 894 86348 900 86351
rect 126 86342 900 86348
rect 1548 86348 1554 86351
rect 1548 86342 1584 86348
rect 126 86308 138 86342
rect 1572 86308 1584 86342
rect 126 86302 900 86308
rect 894 86299 900 86302
rect 1548 86302 1584 86308
rect 1548 86299 1554 86302
rect 156 86262 162 86265
rect 126 86256 162 86262
rect 810 86262 816 86265
rect 810 86256 1584 86262
rect 126 86222 138 86256
rect 1572 86222 1584 86256
rect 126 86216 162 86222
rect 156 86213 162 86216
rect 810 86216 1584 86222
rect 810 86213 816 86216
rect 894 86176 900 86179
rect 126 86170 900 86176
rect 1548 86176 1554 86179
rect 1548 86170 1584 86176
rect 126 86136 138 86170
rect 1572 86136 1584 86170
rect 126 86130 900 86136
rect 894 86127 900 86130
rect 1548 86130 1584 86136
rect 1548 86127 1554 86130
rect 156 86090 162 86093
rect 126 86084 162 86090
rect 810 86090 816 86093
rect 810 86084 1584 86090
rect 126 86050 138 86084
rect 1572 86050 1584 86084
rect 126 86044 162 86050
rect 156 86041 162 86044
rect 810 86044 1584 86050
rect 810 86041 816 86044
rect 894 86004 900 86007
rect 126 85998 900 86004
rect 1548 86004 1554 86007
rect 1548 85998 1584 86004
rect 126 85964 138 85998
rect 1572 85964 1584 85998
rect 126 85958 900 85964
rect 894 85955 900 85958
rect 1548 85958 1584 85964
rect 1548 85955 1554 85958
rect 156 85918 162 85921
rect 126 85912 162 85918
rect 810 85918 816 85921
rect 810 85912 1584 85918
rect 126 85878 138 85912
rect 1572 85878 1584 85912
rect 126 85872 162 85878
rect 156 85869 162 85872
rect 810 85872 1584 85878
rect 810 85869 816 85872
rect 894 85832 900 85835
rect 126 85826 900 85832
rect 1548 85832 1554 85835
rect 1548 85826 1584 85832
rect 126 85792 138 85826
rect 1572 85792 1584 85826
rect 126 85786 900 85792
rect 894 85783 900 85786
rect 1548 85786 1584 85792
rect 1548 85783 1554 85786
rect 156 85746 162 85749
rect 126 85740 162 85746
rect 810 85746 816 85749
rect 810 85740 1584 85746
rect 126 85706 138 85740
rect 1572 85706 1584 85740
rect 126 85700 162 85706
rect 156 85697 162 85700
rect 810 85700 1584 85706
rect 810 85697 816 85700
rect 894 85660 900 85663
rect 126 85654 900 85660
rect 1548 85660 1554 85663
rect 1548 85654 1584 85660
rect 126 85620 138 85654
rect 1572 85620 1584 85654
rect 126 85614 900 85620
rect 894 85611 900 85614
rect 1548 85614 1584 85620
rect 1548 85611 1554 85614
rect 156 85574 162 85577
rect 126 85568 162 85574
rect 810 85574 816 85577
rect 810 85568 1584 85574
rect 126 85534 138 85568
rect 1572 85534 1584 85568
rect 126 85528 162 85534
rect 156 85525 162 85528
rect 810 85528 1584 85534
rect 810 85525 816 85528
rect 894 85488 900 85491
rect 126 85482 900 85488
rect 1548 85488 1554 85491
rect 1548 85482 1584 85488
rect 126 85448 138 85482
rect 1572 85448 1584 85482
rect 126 85442 900 85448
rect 894 85439 900 85442
rect 1548 85442 1584 85448
rect 1548 85439 1554 85442
rect 156 85402 162 85405
rect 126 85396 162 85402
rect 810 85402 816 85405
rect 810 85396 1584 85402
rect 126 85362 138 85396
rect 1572 85362 1584 85396
rect 126 85356 162 85362
rect 156 85353 162 85356
rect 810 85356 1584 85362
rect 810 85353 816 85356
rect 894 85316 900 85319
rect 126 85310 900 85316
rect 1548 85316 1554 85319
rect 1548 85310 1584 85316
rect 126 85276 138 85310
rect 1572 85276 1584 85310
rect 126 85270 900 85276
rect 894 85267 900 85270
rect 1548 85270 1584 85276
rect 1548 85267 1554 85270
rect 156 85230 162 85233
rect 126 85224 162 85230
rect 810 85230 816 85233
rect 810 85224 1584 85230
rect 126 85190 138 85224
rect 1572 85190 1584 85224
rect 126 85184 162 85190
rect 156 85181 162 85184
rect 810 85184 1584 85190
rect 810 85181 816 85184
rect 894 85144 900 85147
rect 126 85138 900 85144
rect 1548 85144 1554 85147
rect 1548 85138 1584 85144
rect 126 85104 138 85138
rect 1572 85104 1584 85138
rect 126 85098 900 85104
rect 894 85095 900 85098
rect 1548 85098 1584 85104
rect 1548 85095 1554 85098
rect 156 85058 162 85061
rect 126 85052 162 85058
rect 810 85058 816 85061
rect 810 85052 1584 85058
rect 126 85018 138 85052
rect 1572 85018 1584 85052
rect 126 85012 162 85018
rect 156 85009 162 85012
rect 810 85012 1584 85018
rect 810 85009 816 85012
rect 894 84972 900 84975
rect 126 84966 900 84972
rect 1548 84972 1554 84975
rect 1548 84966 1584 84972
rect 126 84932 138 84966
rect 1572 84932 1584 84966
rect 126 84926 900 84932
rect 894 84923 900 84926
rect 1548 84926 1584 84932
rect 1548 84923 1554 84926
rect 156 84886 162 84889
rect 126 84880 162 84886
rect 810 84886 816 84889
rect 810 84880 1584 84886
rect 126 84846 138 84880
rect 1572 84846 1584 84880
rect 126 84840 162 84846
rect 156 84837 162 84840
rect 810 84840 1584 84846
rect 810 84837 816 84840
rect 894 84800 900 84803
rect 126 84794 900 84800
rect 1548 84800 1554 84803
rect 1548 84794 1584 84800
rect 126 84760 138 84794
rect 1572 84760 1584 84794
rect 126 84754 900 84760
rect 894 84751 900 84754
rect 1548 84754 1584 84760
rect 1548 84751 1554 84754
rect 156 84714 162 84717
rect 126 84708 162 84714
rect 810 84714 816 84717
rect 810 84708 1584 84714
rect 126 84674 138 84708
rect 1572 84674 1584 84708
rect 126 84668 162 84674
rect 156 84665 162 84668
rect 810 84668 1584 84674
rect 810 84665 816 84668
rect 894 84628 900 84631
rect 126 84622 900 84628
rect 1548 84628 1554 84631
rect 1548 84622 1584 84628
rect 126 84588 138 84622
rect 1572 84588 1584 84622
rect 126 84582 900 84588
rect 894 84579 900 84582
rect 1548 84582 1584 84588
rect 1548 84579 1554 84582
rect 156 84542 162 84545
rect 126 84536 162 84542
rect 810 84542 816 84545
rect 810 84536 1584 84542
rect 126 84502 138 84536
rect 1572 84502 1584 84536
rect 126 84496 162 84502
rect 156 84493 162 84496
rect 810 84496 1584 84502
rect 810 84493 816 84496
rect 894 84456 900 84459
rect 126 84450 900 84456
rect 1548 84456 1554 84459
rect 1548 84450 1584 84456
rect 126 84416 138 84450
rect 1572 84416 1584 84450
rect 126 84410 900 84416
rect 894 84407 900 84410
rect 1548 84410 1584 84416
rect 1548 84407 1554 84410
rect 156 84370 162 84373
rect 126 84364 162 84370
rect 810 84370 816 84373
rect 810 84364 1584 84370
rect 126 84330 138 84364
rect 1572 84330 1584 84364
rect 126 84324 162 84330
rect 156 84321 162 84324
rect 810 84324 1584 84330
rect 810 84321 816 84324
rect 894 84284 900 84287
rect 126 84278 900 84284
rect 1548 84284 1554 84287
rect 1548 84278 1584 84284
rect 126 84244 138 84278
rect 1572 84244 1584 84278
rect 126 84238 900 84244
rect 894 84235 900 84238
rect 1548 84238 1584 84244
rect 1548 84235 1554 84238
rect 156 84198 162 84201
rect 126 84192 162 84198
rect 810 84198 816 84201
rect 810 84192 1584 84198
rect 126 84158 138 84192
rect 1572 84158 1584 84192
rect 126 84152 162 84158
rect 156 84149 162 84152
rect 810 84152 1584 84158
rect 810 84149 816 84152
rect 894 84112 900 84115
rect 126 84106 900 84112
rect 1548 84112 1554 84115
rect 1548 84106 1584 84112
rect 126 84072 138 84106
rect 1572 84072 1584 84106
rect 126 84066 900 84072
rect 894 84063 900 84066
rect 1548 84066 1584 84072
rect 1548 84063 1554 84066
rect 156 84026 162 84029
rect 126 84020 162 84026
rect 810 84026 816 84029
rect 810 84020 1584 84026
rect 126 83986 138 84020
rect 1572 83986 1584 84020
rect 126 83980 162 83986
rect 156 83977 162 83980
rect 810 83980 1584 83986
rect 810 83977 816 83980
rect 894 83940 900 83943
rect 126 83934 900 83940
rect 1548 83940 1554 83943
rect 1548 83934 1584 83940
rect 126 83900 138 83934
rect 1572 83900 1584 83934
rect 126 83894 900 83900
rect 894 83891 900 83894
rect 1548 83894 1584 83900
rect 1548 83891 1554 83894
rect 156 83854 162 83857
rect 126 83848 162 83854
rect 810 83854 816 83857
rect 810 83848 1584 83854
rect 126 83814 138 83848
rect 1572 83814 1584 83848
rect 126 83808 162 83814
rect 156 83805 162 83808
rect 810 83808 1584 83814
rect 810 83805 816 83808
rect 894 83768 900 83771
rect 126 83762 900 83768
rect 1548 83768 1554 83771
rect 1548 83762 1584 83768
rect 126 83728 138 83762
rect 1572 83728 1584 83762
rect 126 83722 900 83728
rect 894 83719 900 83722
rect 1548 83722 1584 83728
rect 1548 83719 1554 83722
rect 156 83682 162 83685
rect 126 83676 162 83682
rect 810 83682 816 83685
rect 810 83676 1584 83682
rect 126 83642 138 83676
rect 1572 83642 1584 83676
rect 126 83636 162 83642
rect 156 83633 162 83636
rect 810 83636 1584 83642
rect 810 83633 816 83636
rect 894 83596 900 83599
rect 126 83590 900 83596
rect 1548 83596 1554 83599
rect 1548 83590 1584 83596
rect 126 83556 138 83590
rect 1572 83556 1584 83590
rect 126 83550 900 83556
rect 894 83547 900 83550
rect 1548 83550 1584 83556
rect 1548 83547 1554 83550
rect 156 83510 162 83513
rect 126 83504 162 83510
rect 810 83510 816 83513
rect 810 83504 1584 83510
rect 126 83470 138 83504
rect 1572 83470 1584 83504
rect 126 83464 162 83470
rect 156 83461 162 83464
rect 810 83464 1584 83470
rect 810 83461 816 83464
rect 894 83424 900 83427
rect 126 83418 900 83424
rect 1548 83424 1554 83427
rect 1548 83418 1584 83424
rect 126 83384 138 83418
rect 1572 83384 1584 83418
rect 126 83378 900 83384
rect 894 83375 900 83378
rect 1548 83378 1584 83384
rect 1548 83375 1554 83378
rect 156 83338 162 83341
rect 126 83332 162 83338
rect 810 83338 816 83341
rect 810 83332 1584 83338
rect 126 83298 138 83332
rect 1572 83298 1584 83332
rect 126 83292 162 83298
rect 156 83289 162 83292
rect 810 83292 1584 83298
rect 810 83289 816 83292
rect 894 83252 900 83255
rect 126 83246 900 83252
rect 1548 83252 1554 83255
rect 1548 83246 1584 83252
rect 126 83212 138 83246
rect 1572 83212 1584 83246
rect 126 83206 900 83212
rect 894 83203 900 83206
rect 1548 83206 1584 83212
rect 1548 83203 1554 83206
rect 156 83166 162 83169
rect 126 83160 162 83166
rect 810 83166 816 83169
rect 810 83160 1584 83166
rect 126 83126 138 83160
rect 1572 83126 1584 83160
rect 126 83120 162 83126
rect 156 83117 162 83120
rect 810 83120 1584 83126
rect 810 83117 816 83120
rect 894 83080 900 83083
rect 126 83074 900 83080
rect 1548 83080 1554 83083
rect 1548 83074 1584 83080
rect 126 83040 138 83074
rect 1572 83040 1584 83074
rect 126 83034 900 83040
rect 894 83031 900 83034
rect 1548 83034 1584 83040
rect 1548 83031 1554 83034
rect 156 82994 162 82997
rect 126 82988 162 82994
rect 810 82994 816 82997
rect 810 82988 1584 82994
rect 126 82954 138 82988
rect 1572 82954 1584 82988
rect 126 82948 162 82954
rect 156 82945 162 82948
rect 810 82948 1584 82954
rect 810 82945 816 82948
rect 894 82908 900 82911
rect 126 82902 900 82908
rect 1548 82908 1554 82911
rect 1548 82902 1584 82908
rect 126 82868 138 82902
rect 1572 82868 1584 82902
rect 126 82862 900 82868
rect 894 82859 900 82862
rect 1548 82862 1584 82868
rect 1548 82859 1554 82862
rect 156 82822 162 82825
rect 126 82816 162 82822
rect 810 82822 816 82825
rect 810 82816 1584 82822
rect 126 82782 138 82816
rect 1572 82782 1584 82816
rect 126 82776 162 82782
rect 156 82773 162 82776
rect 810 82776 1584 82782
rect 810 82773 816 82776
rect 894 82736 900 82739
rect 126 82730 900 82736
rect 1548 82736 1554 82739
rect 1548 82730 1584 82736
rect 126 82696 138 82730
rect 1572 82696 1584 82730
rect 126 82690 900 82696
rect 894 82687 900 82690
rect 1548 82690 1584 82696
rect 1548 82687 1554 82690
rect 156 82650 162 82653
rect 126 82644 162 82650
rect 810 82650 816 82653
rect 810 82644 1584 82650
rect 126 82610 138 82644
rect 1572 82610 1584 82644
rect 126 82604 162 82610
rect 156 82601 162 82604
rect 810 82604 1584 82610
rect 810 82601 816 82604
rect 894 82564 900 82567
rect 126 82558 900 82564
rect 1548 82564 1554 82567
rect 1548 82558 1584 82564
rect 126 82524 138 82558
rect 1572 82524 1584 82558
rect 126 82518 900 82524
rect 894 82515 900 82518
rect 1548 82518 1584 82524
rect 1548 82515 1554 82518
rect 156 82478 162 82481
rect 126 82472 162 82478
rect 810 82478 816 82481
rect 810 82472 1584 82478
rect 126 82438 138 82472
rect 1572 82438 1584 82472
rect 126 82432 162 82438
rect 156 82429 162 82432
rect 810 82432 1584 82438
rect 810 82429 816 82432
rect 894 82392 900 82395
rect 126 82386 900 82392
rect 1548 82392 1554 82395
rect 1548 82386 1584 82392
rect 126 82352 138 82386
rect 1572 82352 1584 82386
rect 126 82346 900 82352
rect 894 82343 900 82346
rect 1548 82346 1584 82352
rect 1548 82343 1554 82346
rect 156 82306 162 82309
rect 126 82300 162 82306
rect 810 82306 816 82309
rect 810 82300 1584 82306
rect 126 82266 138 82300
rect 1572 82266 1584 82300
rect 126 82260 162 82266
rect 156 82257 162 82260
rect 810 82260 1584 82266
rect 810 82257 816 82260
rect 894 82220 900 82223
rect 126 82214 900 82220
rect 1548 82220 1554 82223
rect 1548 82214 1584 82220
rect 126 82180 138 82214
rect 1572 82180 1584 82214
rect 126 82174 900 82180
rect 894 82171 900 82174
rect 1548 82174 1584 82180
rect 1548 82171 1554 82174
rect 156 82134 162 82137
rect 126 82128 162 82134
rect 810 82134 816 82137
rect 810 82128 1584 82134
rect 126 82094 138 82128
rect 1572 82094 1584 82128
rect 126 82088 162 82094
rect 156 82085 162 82088
rect 810 82088 1584 82094
rect 810 82085 816 82088
rect 894 82048 900 82051
rect 126 82042 900 82048
rect 1548 82048 1554 82051
rect 1548 82042 1584 82048
rect 126 82008 138 82042
rect 1572 82008 1584 82042
rect 126 82002 900 82008
rect 894 81999 900 82002
rect 1548 82002 1584 82008
rect 1548 81999 1554 82002
rect 156 81962 162 81965
rect 126 81956 162 81962
rect 810 81962 816 81965
rect 810 81956 1584 81962
rect 126 81922 138 81956
rect 1572 81922 1584 81956
rect 126 81916 162 81922
rect 156 81913 162 81916
rect 810 81916 1584 81922
rect 810 81913 816 81916
rect 894 81876 900 81879
rect 126 81870 900 81876
rect 1548 81876 1554 81879
rect 1548 81870 1584 81876
rect 126 81836 138 81870
rect 1572 81836 1584 81870
rect 126 81830 900 81836
rect 894 81827 900 81830
rect 1548 81830 1584 81836
rect 1548 81827 1554 81830
rect 156 81790 162 81793
rect 126 81784 162 81790
rect 810 81790 816 81793
rect 810 81784 1584 81790
rect 126 81750 138 81784
rect 1572 81750 1584 81784
rect 126 81744 162 81750
rect 156 81741 162 81744
rect 810 81744 1584 81750
rect 810 81741 816 81744
rect 894 81704 900 81707
rect 126 81698 900 81704
rect 1548 81704 1554 81707
rect 1548 81698 1584 81704
rect 126 81664 138 81698
rect 1572 81664 1584 81698
rect 126 81658 900 81664
rect 894 81655 900 81658
rect 1548 81658 1584 81664
rect 1548 81655 1554 81658
rect 156 81618 162 81621
rect 126 81612 162 81618
rect 810 81618 816 81621
rect 810 81612 1584 81618
rect 126 81578 138 81612
rect 1572 81578 1584 81612
rect 126 81572 162 81578
rect 156 81569 162 81572
rect 810 81572 1584 81578
rect 810 81569 816 81572
rect 894 81532 900 81535
rect 126 81526 900 81532
rect 1548 81532 1554 81535
rect 1548 81526 1584 81532
rect 126 81492 138 81526
rect 1572 81492 1584 81526
rect 126 81486 900 81492
rect 894 81483 900 81486
rect 1548 81486 1584 81492
rect 1548 81483 1554 81486
rect 156 81446 162 81449
rect 126 81440 162 81446
rect 810 81446 816 81449
rect 810 81440 1584 81446
rect 126 81406 138 81440
rect 1572 81406 1584 81440
rect 126 81400 162 81406
rect 156 81397 162 81400
rect 810 81400 1584 81406
rect 810 81397 816 81400
rect 894 81360 900 81363
rect 126 81354 900 81360
rect 1548 81360 1554 81363
rect 1548 81354 1584 81360
rect 126 81320 138 81354
rect 1572 81320 1584 81354
rect 126 81314 900 81320
rect 894 81311 900 81314
rect 1548 81314 1584 81320
rect 1548 81311 1554 81314
rect 156 81274 162 81277
rect 126 81268 162 81274
rect 810 81274 816 81277
rect 810 81268 1584 81274
rect 126 81234 138 81268
rect 1572 81234 1584 81268
rect 126 81228 162 81234
rect 156 81225 162 81228
rect 810 81228 1584 81234
rect 810 81225 816 81228
rect 894 81188 900 81191
rect 126 81182 900 81188
rect 1548 81188 1554 81191
rect 1548 81182 1584 81188
rect 126 81148 138 81182
rect 1572 81148 1584 81182
rect 126 81142 900 81148
rect 894 81139 900 81142
rect 1548 81142 1584 81148
rect 1548 81139 1554 81142
rect 156 81102 162 81105
rect 126 81096 162 81102
rect 810 81102 816 81105
rect 810 81096 1584 81102
rect 126 81062 138 81096
rect 1572 81062 1584 81096
rect 126 81056 162 81062
rect 156 81053 162 81056
rect 810 81056 1584 81062
rect 810 81053 816 81056
rect 894 81016 900 81019
rect 126 81010 900 81016
rect 1548 81016 1554 81019
rect 1548 81010 1584 81016
rect 126 80976 138 81010
rect 1572 80976 1584 81010
rect 126 80970 900 80976
rect 894 80967 900 80970
rect 1548 80970 1584 80976
rect 1548 80967 1554 80970
rect 156 80930 162 80933
rect 126 80924 162 80930
rect 810 80930 816 80933
rect 810 80924 1584 80930
rect 126 80890 138 80924
rect 1572 80890 1584 80924
rect 126 80884 162 80890
rect 156 80881 162 80884
rect 810 80884 1584 80890
rect 810 80881 816 80884
rect 894 80844 900 80847
rect 126 80838 900 80844
rect 1548 80844 1554 80847
rect 1548 80838 1584 80844
rect 126 80804 138 80838
rect 1572 80804 1584 80838
rect 126 80798 900 80804
rect 894 80795 900 80798
rect 1548 80798 1584 80804
rect 1548 80795 1554 80798
rect 156 80758 162 80761
rect 126 80752 162 80758
rect 810 80758 816 80761
rect 810 80752 1584 80758
rect 126 80718 138 80752
rect 1572 80718 1584 80752
rect 126 80712 162 80718
rect 156 80709 162 80712
rect 810 80712 1584 80718
rect 810 80709 816 80712
rect 894 80672 900 80675
rect 126 80666 900 80672
rect 1548 80672 1554 80675
rect 1548 80666 1584 80672
rect 126 80632 138 80666
rect 1572 80632 1584 80666
rect 126 80626 900 80632
rect 894 80623 900 80626
rect 1548 80626 1584 80632
rect 1548 80623 1554 80626
rect 156 80586 162 80589
rect 126 80580 162 80586
rect 810 80586 816 80589
rect 810 80580 1584 80586
rect 126 80546 138 80580
rect 1572 80546 1584 80580
rect 126 80540 162 80546
rect 156 80537 162 80540
rect 810 80540 1584 80546
rect 810 80537 816 80540
rect 894 80500 900 80503
rect 126 80494 900 80500
rect 1548 80500 1554 80503
rect 1548 80494 1584 80500
rect 126 80460 138 80494
rect 1572 80460 1584 80494
rect 126 80454 900 80460
rect 894 80451 900 80454
rect 1548 80454 1584 80460
rect 1548 80451 1554 80454
rect 156 80414 162 80417
rect 126 80408 162 80414
rect 810 80414 816 80417
rect 810 80408 1584 80414
rect 126 80374 138 80408
rect 1572 80374 1584 80408
rect 126 80368 162 80374
rect 156 80365 162 80368
rect 810 80368 1584 80374
rect 810 80365 816 80368
rect 894 80328 900 80331
rect 126 80322 900 80328
rect 1548 80328 1554 80331
rect 1548 80322 1584 80328
rect 126 80288 138 80322
rect 1572 80288 1584 80322
rect 126 80282 900 80288
rect 894 80279 900 80282
rect 1548 80282 1584 80288
rect 1548 80279 1554 80282
rect 156 80242 162 80245
rect 126 80236 162 80242
rect 810 80242 816 80245
rect 810 80236 1584 80242
rect 126 80202 138 80236
rect 1572 80202 1584 80236
rect 126 80196 162 80202
rect 156 80193 162 80196
rect 810 80196 1584 80202
rect 810 80193 816 80196
rect 894 80156 900 80159
rect 126 80150 900 80156
rect 1548 80156 1554 80159
rect 1548 80150 1584 80156
rect 126 80116 138 80150
rect 1572 80116 1584 80150
rect 126 80110 900 80116
rect 894 80107 900 80110
rect 1548 80110 1584 80116
rect 1548 80107 1554 80110
rect 156 80070 162 80073
rect 126 80064 162 80070
rect 810 80070 816 80073
rect 810 80064 1584 80070
rect 126 80030 138 80064
rect 1572 80030 1584 80064
rect 126 80024 162 80030
rect 156 80021 162 80024
rect 810 80024 1584 80030
rect 810 80021 816 80024
rect 894 79984 900 79987
rect 126 79978 900 79984
rect 1548 79984 1554 79987
rect 1548 79978 1584 79984
rect 126 79944 138 79978
rect 1572 79944 1584 79978
rect 126 79938 900 79944
rect 894 79935 900 79938
rect 1548 79938 1584 79944
rect 1548 79935 1554 79938
rect 156 79898 162 79901
rect 126 79892 162 79898
rect 810 79898 816 79901
rect 810 79892 1584 79898
rect 126 79858 138 79892
rect 1572 79858 1584 79892
rect 126 79852 162 79858
rect 156 79849 162 79852
rect 810 79852 1584 79858
rect 810 79849 816 79852
rect 894 79812 900 79815
rect 126 79806 900 79812
rect 1548 79812 1554 79815
rect 1548 79806 1584 79812
rect 126 79772 138 79806
rect 1572 79772 1584 79806
rect 126 79766 900 79772
rect 894 79763 900 79766
rect 1548 79766 1584 79772
rect 1548 79763 1554 79766
rect 156 79726 162 79729
rect 126 79720 162 79726
rect 810 79726 816 79729
rect 810 79720 1584 79726
rect 126 79686 138 79720
rect 1572 79686 1584 79720
rect 126 79680 162 79686
rect 156 79677 162 79680
rect 810 79680 1584 79686
rect 810 79677 816 79680
rect 894 79640 900 79643
rect 126 79634 900 79640
rect 1548 79640 1554 79643
rect 1548 79634 1584 79640
rect 126 79600 138 79634
rect 1572 79600 1584 79634
rect 126 79594 900 79600
rect 894 79591 900 79594
rect 1548 79594 1584 79600
rect 1548 79591 1554 79594
rect 156 79554 162 79557
rect 126 79548 162 79554
rect 810 79554 816 79557
rect 810 79548 1584 79554
rect 126 79514 138 79548
rect 1572 79514 1584 79548
rect 126 79508 162 79514
rect 156 79505 162 79508
rect 810 79508 1584 79514
rect 810 79505 816 79508
rect 894 79468 900 79471
rect 126 79462 900 79468
rect 1548 79468 1554 79471
rect 1548 79462 1584 79468
rect 126 79428 138 79462
rect 1572 79428 1584 79462
rect 126 79422 900 79428
rect 894 79419 900 79422
rect 1548 79422 1584 79428
rect 1548 79419 1554 79422
rect 156 79382 162 79385
rect 126 79376 162 79382
rect 810 79382 816 79385
rect 810 79376 1584 79382
rect 126 79342 138 79376
rect 1572 79342 1584 79376
rect 126 79336 162 79342
rect 156 79333 162 79336
rect 810 79336 1584 79342
rect 810 79333 816 79336
rect 894 79296 900 79299
rect 126 79290 900 79296
rect 1548 79296 1554 79299
rect 1548 79290 1584 79296
rect 126 79256 138 79290
rect 1572 79256 1584 79290
rect 126 79250 900 79256
rect 894 79247 900 79250
rect 1548 79250 1584 79256
rect 1548 79247 1554 79250
rect 156 79210 162 79213
rect 126 79204 162 79210
rect 810 79210 816 79213
rect 810 79204 1584 79210
rect 126 79170 138 79204
rect 1572 79170 1584 79204
rect 126 79164 162 79170
rect 156 79161 162 79164
rect 810 79164 1584 79170
rect 810 79161 816 79164
rect 894 79124 900 79127
rect 126 79118 900 79124
rect 1548 79124 1554 79127
rect 1548 79118 1584 79124
rect 126 79084 138 79118
rect 1572 79084 1584 79118
rect 126 79078 900 79084
rect 894 79075 900 79078
rect 1548 79078 1584 79084
rect 1548 79075 1554 79078
rect 156 79038 162 79041
rect 126 79032 162 79038
rect 810 79038 816 79041
rect 810 79032 1584 79038
rect 126 78998 138 79032
rect 1572 78998 1584 79032
rect 126 78992 162 78998
rect 156 78989 162 78992
rect 810 78992 1584 78998
rect 810 78989 816 78992
rect 894 78952 900 78955
rect 126 78946 900 78952
rect 1548 78952 1554 78955
rect 1548 78946 1584 78952
rect 126 78912 138 78946
rect 1572 78912 1584 78946
rect 126 78906 900 78912
rect 894 78903 900 78906
rect 1548 78906 1584 78912
rect 1548 78903 1554 78906
rect 156 78866 162 78869
rect 126 78860 162 78866
rect 810 78866 816 78869
rect 810 78860 1584 78866
rect 126 78826 138 78860
rect 1572 78826 1584 78860
rect 126 78820 162 78826
rect 156 78817 162 78820
rect 810 78820 1584 78826
rect 810 78817 816 78820
rect 894 78780 900 78783
rect 126 78774 900 78780
rect 1548 78780 1554 78783
rect 1548 78774 1584 78780
rect 126 78740 138 78774
rect 1572 78740 1584 78774
rect 126 78734 900 78740
rect 894 78731 900 78734
rect 1548 78734 1584 78740
rect 1548 78731 1554 78734
rect 156 78694 162 78697
rect 126 78688 162 78694
rect 810 78694 816 78697
rect 810 78688 1584 78694
rect 126 78654 138 78688
rect 1572 78654 1584 78688
rect 126 78648 162 78654
rect 156 78645 162 78648
rect 810 78648 1584 78654
rect 810 78645 816 78648
rect 894 78608 900 78611
rect 126 78602 900 78608
rect 1548 78608 1554 78611
rect 1548 78602 1584 78608
rect 126 78568 138 78602
rect 1572 78568 1584 78602
rect 126 78562 900 78568
rect 894 78559 900 78562
rect 1548 78562 1584 78568
rect 1548 78559 1554 78562
rect 156 78522 162 78525
rect 126 78516 162 78522
rect 810 78522 816 78525
rect 810 78516 1584 78522
rect 126 78482 138 78516
rect 1572 78482 1584 78516
rect 126 78476 162 78482
rect 156 78473 162 78476
rect 810 78476 1584 78482
rect 810 78473 816 78476
rect 894 78436 900 78439
rect 126 78430 900 78436
rect 1548 78436 1554 78439
rect 1548 78430 1584 78436
rect 126 78396 138 78430
rect 1572 78396 1584 78430
rect 126 78390 900 78396
rect 894 78387 900 78390
rect 1548 78390 1584 78396
rect 1548 78387 1554 78390
rect 156 78350 162 78353
rect 126 78344 162 78350
rect 810 78350 816 78353
rect 810 78344 1584 78350
rect 126 78310 138 78344
rect 1572 78310 1584 78344
rect 126 78304 162 78310
rect 156 78301 162 78304
rect 810 78304 1584 78310
rect 810 78301 816 78304
rect 894 78264 900 78267
rect 126 78258 900 78264
rect 1548 78264 1554 78267
rect 1548 78258 1584 78264
rect 126 78224 138 78258
rect 1572 78224 1584 78258
rect 126 78218 900 78224
rect 894 78215 900 78218
rect 1548 78218 1584 78224
rect 1548 78215 1554 78218
rect 156 78178 162 78181
rect 126 78172 162 78178
rect 810 78178 816 78181
rect 810 78172 1584 78178
rect 126 78138 138 78172
rect 1572 78138 1584 78172
rect 126 78132 162 78138
rect 156 78129 162 78132
rect 810 78132 1584 78138
rect 810 78129 816 78132
rect 894 78092 900 78095
rect 126 78086 900 78092
rect 1548 78092 1554 78095
rect 1548 78086 1584 78092
rect 126 78052 138 78086
rect 1572 78052 1584 78086
rect 126 78046 900 78052
rect 894 78043 900 78046
rect 1548 78046 1584 78052
rect 1548 78043 1554 78046
rect 156 78006 162 78009
rect 126 78000 162 78006
rect 810 78006 816 78009
rect 810 78000 1584 78006
rect 126 77966 138 78000
rect 1572 77966 1584 78000
rect 126 77960 162 77966
rect 156 77957 162 77960
rect 810 77960 1584 77966
rect 810 77957 816 77960
rect 894 77920 900 77923
rect 126 77914 900 77920
rect 1548 77920 1554 77923
rect 1548 77914 1584 77920
rect 126 77880 138 77914
rect 1572 77880 1584 77914
rect 126 77874 900 77880
rect 894 77871 900 77874
rect 1548 77874 1584 77880
rect 1548 77871 1554 77874
rect 156 77834 162 77837
rect 126 77828 162 77834
rect 810 77834 816 77837
rect 810 77828 1584 77834
rect 126 77794 138 77828
rect 1572 77794 1584 77828
rect 126 77788 162 77794
rect 156 77785 162 77788
rect 810 77788 1584 77794
rect 810 77785 816 77788
rect 894 77748 900 77751
rect 126 77742 900 77748
rect 1548 77748 1554 77751
rect 1548 77742 1584 77748
rect 126 77708 138 77742
rect 1572 77708 1584 77742
rect 126 77702 900 77708
rect 894 77699 900 77702
rect 1548 77702 1584 77708
rect 1548 77699 1554 77702
rect 156 77662 162 77665
rect 126 77656 162 77662
rect 810 77662 816 77665
rect 810 77656 1584 77662
rect 126 77622 138 77656
rect 1572 77622 1584 77656
rect 126 77616 162 77622
rect 156 77613 162 77616
rect 810 77616 1584 77622
rect 810 77613 816 77616
rect 894 77576 900 77579
rect 126 77570 900 77576
rect 1548 77576 1554 77579
rect 1548 77570 1584 77576
rect 126 77536 138 77570
rect 1572 77536 1584 77570
rect 126 77530 900 77536
rect 894 77527 900 77530
rect 1548 77530 1584 77536
rect 1548 77527 1554 77530
rect 156 77490 162 77493
rect 126 77484 162 77490
rect 810 77490 816 77493
rect 810 77484 1584 77490
rect 126 77450 138 77484
rect 1572 77450 1584 77484
rect 126 77444 162 77450
rect 156 77441 162 77444
rect 810 77444 1584 77450
rect 810 77441 816 77444
rect 894 77404 900 77407
rect 126 77398 900 77404
rect 1548 77404 1554 77407
rect 1548 77398 1584 77404
rect 126 77364 138 77398
rect 1572 77364 1584 77398
rect 126 77358 900 77364
rect 894 77355 900 77358
rect 1548 77358 1584 77364
rect 1548 77355 1554 77358
rect 156 77318 162 77321
rect 126 77312 162 77318
rect 810 77318 816 77321
rect 810 77312 1584 77318
rect 126 77278 138 77312
rect 1572 77278 1584 77312
rect 126 77272 162 77278
rect 156 77269 162 77272
rect 810 77272 1584 77278
rect 810 77269 816 77272
rect 894 77232 900 77235
rect 126 77226 900 77232
rect 1548 77232 1554 77235
rect 1548 77226 1584 77232
rect 126 77192 138 77226
rect 1572 77192 1584 77226
rect 126 77186 900 77192
rect 894 77183 900 77186
rect 1548 77186 1584 77192
rect 1548 77183 1554 77186
rect 156 77146 162 77149
rect 126 77140 162 77146
rect 810 77146 816 77149
rect 810 77140 1584 77146
rect 126 77106 138 77140
rect 1572 77106 1584 77140
rect 126 77100 162 77106
rect 156 77097 162 77100
rect 810 77100 1584 77106
rect 810 77097 816 77100
rect 894 77060 900 77063
rect 126 77054 900 77060
rect 1548 77060 1554 77063
rect 1548 77054 1584 77060
rect 126 77020 138 77054
rect 1572 77020 1584 77054
rect 126 77014 900 77020
rect 894 77011 900 77014
rect 1548 77014 1584 77020
rect 1548 77011 1554 77014
rect 156 76974 162 76977
rect 126 76968 162 76974
rect 810 76974 816 76977
rect 810 76968 1584 76974
rect 126 76934 138 76968
rect 1572 76934 1584 76968
rect 126 76928 162 76934
rect 156 76925 162 76928
rect 810 76928 1584 76934
rect 810 76925 816 76928
rect 894 76888 900 76891
rect 126 76882 900 76888
rect 1548 76888 1554 76891
rect 1548 76882 1584 76888
rect 126 76848 138 76882
rect 1572 76848 1584 76882
rect 126 76842 900 76848
rect 894 76839 900 76842
rect 1548 76842 1584 76848
rect 1548 76839 1554 76842
rect 156 76802 162 76805
rect 126 76796 162 76802
rect 810 76802 816 76805
rect 810 76796 1584 76802
rect 126 76762 138 76796
rect 1572 76762 1584 76796
rect 126 76756 162 76762
rect 156 76753 162 76756
rect 810 76756 1584 76762
rect 810 76753 816 76756
rect 894 76716 900 76719
rect 126 76710 900 76716
rect 1548 76716 1554 76719
rect 1548 76710 1584 76716
rect 126 76676 138 76710
rect 1572 76676 1584 76710
rect 126 76670 900 76676
rect 894 76667 900 76670
rect 1548 76670 1584 76676
rect 1548 76667 1554 76670
rect 156 76630 162 76633
rect 126 76624 162 76630
rect 810 76630 816 76633
rect 810 76624 1584 76630
rect 126 76590 138 76624
rect 1572 76590 1584 76624
rect 126 76584 162 76590
rect 156 76581 162 76584
rect 810 76584 1584 76590
rect 810 76581 816 76584
rect 894 76544 900 76547
rect 126 76538 900 76544
rect 1548 76544 1554 76547
rect 1548 76538 1584 76544
rect 126 76504 138 76538
rect 1572 76504 1584 76538
rect 126 76498 900 76504
rect 894 76495 900 76498
rect 1548 76498 1584 76504
rect 1548 76495 1554 76498
rect 156 76458 162 76461
rect 126 76452 162 76458
rect 810 76458 816 76461
rect 810 76452 1584 76458
rect 126 76418 138 76452
rect 1572 76418 1584 76452
rect 126 76412 162 76418
rect 156 76409 162 76412
rect 810 76412 1584 76418
rect 810 76409 816 76412
rect 894 76372 900 76375
rect 126 76366 900 76372
rect 1548 76372 1554 76375
rect 1548 76366 1584 76372
rect 126 76332 138 76366
rect 1572 76332 1584 76366
rect 126 76326 900 76332
rect 894 76323 900 76326
rect 1548 76326 1584 76332
rect 1548 76323 1554 76326
rect 156 76286 162 76289
rect 126 76280 162 76286
rect 810 76286 816 76289
rect 810 76280 1584 76286
rect 126 76246 138 76280
rect 1572 76246 1584 76280
rect 126 76240 162 76246
rect 156 76237 162 76240
rect 810 76240 1584 76246
rect 810 76237 816 76240
rect 894 76200 900 76203
rect 126 76194 900 76200
rect 1548 76200 1554 76203
rect 1548 76194 1584 76200
rect 126 76160 138 76194
rect 1572 76160 1584 76194
rect 126 76154 900 76160
rect 894 76151 900 76154
rect 1548 76154 1584 76160
rect 1548 76151 1554 76154
rect 156 76114 162 76117
rect 126 76108 162 76114
rect 810 76114 816 76117
rect 810 76108 1584 76114
rect 126 76074 138 76108
rect 1572 76074 1584 76108
rect 126 76068 162 76074
rect 156 76065 162 76068
rect 810 76068 1584 76074
rect 810 76065 816 76068
rect 894 76028 900 76031
rect 126 76022 900 76028
rect 1548 76028 1554 76031
rect 1548 76022 1584 76028
rect 126 75988 138 76022
rect 1572 75988 1584 76022
rect 126 75982 900 75988
rect 894 75979 900 75982
rect 1548 75982 1584 75988
rect 1548 75979 1554 75982
rect 156 75942 162 75945
rect 126 75936 162 75942
rect 810 75942 816 75945
rect 810 75936 1584 75942
rect 126 75902 138 75936
rect 1572 75902 1584 75936
rect 126 75896 162 75902
rect 156 75893 162 75896
rect 810 75896 1584 75902
rect 810 75893 816 75896
rect 894 75856 900 75859
rect 126 75850 900 75856
rect 1548 75856 1554 75859
rect 1548 75850 1584 75856
rect 126 75816 138 75850
rect 1572 75816 1584 75850
rect 126 75810 900 75816
rect 894 75807 900 75810
rect 1548 75810 1584 75816
rect 1548 75807 1554 75810
rect 156 75770 162 75773
rect 126 75764 162 75770
rect 810 75770 816 75773
rect 810 75764 1584 75770
rect 126 75730 138 75764
rect 1572 75730 1584 75764
rect 126 75724 162 75730
rect 156 75721 162 75724
rect 810 75724 1584 75730
rect 810 75721 816 75724
rect 894 75684 900 75687
rect 126 75678 900 75684
rect 1548 75684 1554 75687
rect 1548 75678 1584 75684
rect 126 75644 138 75678
rect 1572 75644 1584 75678
rect 126 75638 900 75644
rect 894 75635 900 75638
rect 1548 75638 1584 75644
rect 1548 75635 1554 75638
rect 156 75598 162 75601
rect 126 75592 162 75598
rect 810 75598 816 75601
rect 810 75592 1584 75598
rect 126 75558 138 75592
rect 1572 75558 1584 75592
rect 126 75552 162 75558
rect 156 75549 162 75552
rect 810 75552 1584 75558
rect 810 75549 816 75552
rect 894 75512 900 75515
rect 126 75506 900 75512
rect 1548 75512 1554 75515
rect 1548 75506 1584 75512
rect 126 75472 138 75506
rect 1572 75472 1584 75506
rect 126 75466 900 75472
rect 894 75463 900 75466
rect 1548 75466 1584 75472
rect 1548 75463 1554 75466
rect 156 75426 162 75429
rect 126 75420 162 75426
rect 810 75426 816 75429
rect 810 75420 1584 75426
rect 126 75386 138 75420
rect 1572 75386 1584 75420
rect 126 75380 162 75386
rect 156 75377 162 75380
rect 810 75380 1584 75386
rect 810 75377 816 75380
rect 894 75340 900 75343
rect 126 75334 900 75340
rect 1548 75340 1554 75343
rect 1548 75334 1584 75340
rect 126 75300 138 75334
rect 1572 75300 1584 75334
rect 126 75294 900 75300
rect 894 75291 900 75294
rect 1548 75294 1584 75300
rect 1548 75291 1554 75294
rect 156 75254 162 75257
rect 126 75248 162 75254
rect 810 75254 816 75257
rect 810 75248 1584 75254
rect 126 75214 138 75248
rect 1572 75214 1584 75248
rect 126 75208 162 75214
rect 156 75205 162 75208
rect 810 75208 1584 75214
rect 810 75205 816 75208
rect 894 75168 900 75171
rect 126 75162 900 75168
rect 1548 75168 1554 75171
rect 1548 75162 1584 75168
rect 126 75128 138 75162
rect 1572 75128 1584 75162
rect 126 75122 900 75128
rect 894 75119 900 75122
rect 1548 75122 1584 75128
rect 1548 75119 1554 75122
rect 156 75082 162 75085
rect 126 75076 162 75082
rect 810 75082 816 75085
rect 810 75076 1584 75082
rect 126 75042 138 75076
rect 1572 75042 1584 75076
rect 126 75036 162 75042
rect 156 75033 162 75036
rect 810 75036 1584 75042
rect 810 75033 816 75036
rect 894 74996 900 74999
rect 126 74990 900 74996
rect 1548 74996 1554 74999
rect 1548 74990 1584 74996
rect 126 74956 138 74990
rect 1572 74956 1584 74990
rect 126 74950 900 74956
rect 894 74947 900 74950
rect 1548 74950 1584 74956
rect 1548 74947 1554 74950
rect 156 74910 162 74913
rect 126 74904 162 74910
rect 810 74910 816 74913
rect 810 74904 1584 74910
rect 126 74870 138 74904
rect 1572 74870 1584 74904
rect 126 74864 162 74870
rect 156 74861 162 74864
rect 810 74864 1584 74870
rect 810 74861 816 74864
rect 894 74824 900 74827
rect 126 74818 900 74824
rect 1548 74824 1554 74827
rect 1548 74818 1584 74824
rect 126 74784 138 74818
rect 1572 74784 1584 74818
rect 126 74778 900 74784
rect 894 74775 900 74778
rect 1548 74778 1584 74784
rect 1548 74775 1554 74778
rect 156 74738 162 74741
rect 126 74732 162 74738
rect 810 74738 816 74741
rect 810 74732 1584 74738
rect 126 74698 138 74732
rect 1572 74698 1584 74732
rect 126 74692 162 74698
rect 156 74689 162 74692
rect 810 74692 1584 74698
rect 810 74689 816 74692
rect 894 74652 900 74655
rect 126 74646 900 74652
rect 1548 74652 1554 74655
rect 1548 74646 1584 74652
rect 126 74612 138 74646
rect 1572 74612 1584 74646
rect 126 74606 900 74612
rect 894 74603 900 74606
rect 1548 74606 1584 74612
rect 1548 74603 1554 74606
rect 156 74566 162 74569
rect 126 74560 162 74566
rect 810 74566 816 74569
rect 810 74560 1584 74566
rect 126 74526 138 74560
rect 1572 74526 1584 74560
rect 126 74520 162 74526
rect 156 74517 162 74520
rect 810 74520 1584 74526
rect 810 74517 816 74520
rect 894 74480 900 74483
rect 126 74474 900 74480
rect 1548 74480 1554 74483
rect 1548 74474 1584 74480
rect 126 74440 138 74474
rect 1572 74440 1584 74474
rect 126 74434 900 74440
rect 894 74431 900 74434
rect 1548 74434 1584 74440
rect 1548 74431 1554 74434
rect 156 74394 162 74397
rect 126 74388 162 74394
rect 810 74394 816 74397
rect 810 74388 1584 74394
rect 126 74354 138 74388
rect 1572 74354 1584 74388
rect 126 74348 162 74354
rect 156 74345 162 74348
rect 810 74348 1584 74354
rect 810 74345 816 74348
rect 894 74308 900 74311
rect 126 74302 900 74308
rect 1548 74308 1554 74311
rect 1548 74302 1584 74308
rect 126 74268 138 74302
rect 1572 74268 1584 74302
rect 126 74262 900 74268
rect 894 74259 900 74262
rect 1548 74262 1584 74268
rect 1548 74259 1554 74262
rect 156 74222 162 74225
rect 126 74216 162 74222
rect 810 74222 816 74225
rect 810 74216 1584 74222
rect 126 74182 138 74216
rect 1572 74182 1584 74216
rect 126 74176 162 74182
rect 156 74173 162 74176
rect 810 74176 1584 74182
rect 810 74173 816 74176
rect 894 74136 900 74139
rect 126 74130 900 74136
rect 1548 74136 1554 74139
rect 1548 74130 1584 74136
rect 126 74096 138 74130
rect 1572 74096 1584 74130
rect 126 74090 900 74096
rect 894 74087 900 74090
rect 1548 74090 1584 74096
rect 1548 74087 1554 74090
rect 156 74050 162 74053
rect 126 74044 162 74050
rect 810 74050 816 74053
rect 810 74044 1584 74050
rect 126 74010 138 74044
rect 1572 74010 1584 74044
rect 126 74004 162 74010
rect 156 74001 162 74004
rect 810 74004 1584 74010
rect 810 74001 816 74004
rect 894 73964 900 73967
rect 126 73958 900 73964
rect 1548 73964 1554 73967
rect 1548 73958 1584 73964
rect 126 73924 138 73958
rect 1572 73924 1584 73958
rect 126 73918 900 73924
rect 894 73915 900 73918
rect 1548 73918 1584 73924
rect 1548 73915 1554 73918
rect 156 73878 162 73881
rect 126 73872 162 73878
rect 810 73878 816 73881
rect 810 73872 1584 73878
rect 126 73838 138 73872
rect 1572 73838 1584 73872
rect 126 73832 162 73838
rect 156 73829 162 73832
rect 810 73832 1584 73838
rect 810 73829 816 73832
rect 894 73792 900 73795
rect 126 73786 900 73792
rect 1548 73792 1554 73795
rect 1548 73786 1584 73792
rect 126 73752 138 73786
rect 1572 73752 1584 73786
rect 126 73746 900 73752
rect 894 73743 900 73746
rect 1548 73746 1584 73752
rect 1548 73743 1554 73746
rect 156 73706 162 73709
rect 126 73700 162 73706
rect 810 73706 816 73709
rect 810 73700 1584 73706
rect 126 73666 138 73700
rect 1572 73666 1584 73700
rect 126 73660 162 73666
rect 156 73657 162 73660
rect 810 73660 1584 73666
rect 810 73657 816 73660
rect 894 73620 900 73623
rect 126 73614 900 73620
rect 1548 73620 1554 73623
rect 1548 73614 1584 73620
rect 126 73580 138 73614
rect 1572 73580 1584 73614
rect 126 73574 900 73580
rect 894 73571 900 73574
rect 1548 73574 1584 73580
rect 1548 73571 1554 73574
rect 156 73534 162 73537
rect 126 73528 162 73534
rect 810 73534 816 73537
rect 810 73528 1584 73534
rect 126 73494 138 73528
rect 1572 73494 1584 73528
rect 126 73488 162 73494
rect 156 73485 162 73488
rect 810 73488 1584 73494
rect 810 73485 816 73488
rect 894 73448 900 73451
rect 126 73442 900 73448
rect 1548 73448 1554 73451
rect 1548 73442 1584 73448
rect 126 73408 138 73442
rect 1572 73408 1584 73442
rect 126 73402 900 73408
rect 894 73399 900 73402
rect 1548 73402 1584 73408
rect 1548 73399 1554 73402
rect 156 73362 162 73365
rect 126 73356 162 73362
rect 810 73362 816 73365
rect 810 73356 1584 73362
rect 126 73322 138 73356
rect 1572 73322 1584 73356
rect 126 73316 162 73322
rect 156 73313 162 73316
rect 810 73316 1584 73322
rect 810 73313 816 73316
rect 894 73276 900 73279
rect 126 73270 900 73276
rect 1548 73276 1554 73279
rect 1548 73270 1584 73276
rect 126 73236 138 73270
rect 1572 73236 1584 73270
rect 126 73230 900 73236
rect 894 73227 900 73230
rect 1548 73230 1584 73236
rect 1548 73227 1554 73230
rect 156 73190 162 73193
rect 126 73184 162 73190
rect 810 73190 816 73193
rect 810 73184 1584 73190
rect 126 73150 138 73184
rect 1572 73150 1584 73184
rect 126 73144 162 73150
rect 156 73141 162 73144
rect 810 73144 1584 73150
rect 810 73141 816 73144
rect 894 73104 900 73107
rect 126 73098 900 73104
rect 1548 73104 1554 73107
rect 1548 73098 1584 73104
rect 126 73064 138 73098
rect 1572 73064 1584 73098
rect 126 73058 900 73064
rect 894 73055 900 73058
rect 1548 73058 1584 73064
rect 1548 73055 1554 73058
rect 156 73018 162 73021
rect 126 73012 162 73018
rect 810 73018 816 73021
rect 810 73012 1584 73018
rect 126 72978 138 73012
rect 1572 72978 1584 73012
rect 126 72972 162 72978
rect 156 72969 162 72972
rect 810 72972 1584 72978
rect 810 72969 816 72972
rect 894 72932 900 72935
rect 126 72926 900 72932
rect 1548 72932 1554 72935
rect 1548 72926 1584 72932
rect 126 72892 138 72926
rect 1572 72892 1584 72926
rect 126 72886 900 72892
rect 894 72883 900 72886
rect 1548 72886 1584 72892
rect 1548 72883 1554 72886
rect 156 72846 162 72849
rect 126 72840 162 72846
rect 810 72846 816 72849
rect 810 72840 1584 72846
rect 126 72806 138 72840
rect 1572 72806 1584 72840
rect 126 72800 162 72806
rect 156 72797 162 72800
rect 810 72800 1584 72806
rect 810 72797 816 72800
rect 894 72760 900 72763
rect 126 72754 900 72760
rect 1548 72760 1554 72763
rect 1548 72754 1584 72760
rect 126 72720 138 72754
rect 1572 72720 1584 72754
rect 126 72714 900 72720
rect 894 72711 900 72714
rect 1548 72714 1584 72720
rect 1548 72711 1554 72714
rect 156 72674 162 72677
rect 126 72668 162 72674
rect 810 72674 816 72677
rect 810 72668 1584 72674
rect 126 72634 138 72668
rect 1572 72634 1584 72668
rect 126 72628 162 72634
rect 156 72625 162 72628
rect 810 72628 1584 72634
rect 810 72625 816 72628
rect 894 72588 900 72591
rect 126 72582 900 72588
rect 1548 72588 1554 72591
rect 1548 72582 1584 72588
rect 126 72548 138 72582
rect 1572 72548 1584 72582
rect 126 72542 900 72548
rect 894 72539 900 72542
rect 1548 72542 1584 72548
rect 1548 72539 1554 72542
rect 156 72502 162 72505
rect 126 72496 162 72502
rect 810 72502 816 72505
rect 810 72496 1584 72502
rect 126 72462 138 72496
rect 1572 72462 1584 72496
rect 126 72456 162 72462
rect 156 72453 162 72456
rect 810 72456 1584 72462
rect 810 72453 816 72456
rect 894 72416 900 72419
rect 126 72410 900 72416
rect 1548 72416 1554 72419
rect 1548 72410 1584 72416
rect 126 72376 138 72410
rect 1572 72376 1584 72410
rect 126 72370 900 72376
rect 894 72367 900 72370
rect 1548 72370 1584 72376
rect 1548 72367 1554 72370
rect 156 72330 162 72333
rect 126 72324 162 72330
rect 810 72330 816 72333
rect 810 72324 1584 72330
rect 126 72290 138 72324
rect 1572 72290 1584 72324
rect 126 72284 162 72290
rect 156 72281 162 72284
rect 810 72284 1584 72290
rect 810 72281 816 72284
rect 894 72244 900 72247
rect 126 72238 900 72244
rect 1548 72244 1554 72247
rect 1548 72238 1584 72244
rect 126 72204 138 72238
rect 1572 72204 1584 72238
rect 126 72198 900 72204
rect 894 72195 900 72198
rect 1548 72198 1584 72204
rect 1548 72195 1554 72198
rect 156 72158 162 72161
rect 126 72152 162 72158
rect 810 72158 816 72161
rect 810 72152 1584 72158
rect 126 72118 138 72152
rect 1572 72118 1584 72152
rect 126 72112 162 72118
rect 156 72109 162 72112
rect 810 72112 1584 72118
rect 810 72109 816 72112
rect 894 72072 900 72075
rect 126 72066 900 72072
rect 1548 72072 1554 72075
rect 1548 72066 1584 72072
rect 126 72032 138 72066
rect 1572 72032 1584 72066
rect 126 72026 900 72032
rect 894 72023 900 72026
rect 1548 72026 1584 72032
rect 1548 72023 1554 72026
rect 156 71986 162 71989
rect 126 71980 162 71986
rect 810 71986 816 71989
rect 810 71980 1584 71986
rect 126 71946 138 71980
rect 1572 71946 1584 71980
rect 126 71940 162 71946
rect 156 71937 162 71940
rect 810 71940 1584 71946
rect 810 71937 816 71940
rect 894 71900 900 71903
rect 126 71894 900 71900
rect 1548 71900 1554 71903
rect 1548 71894 1584 71900
rect 126 71860 138 71894
rect 1572 71860 1584 71894
rect 126 71854 900 71860
rect 894 71851 900 71854
rect 1548 71854 1584 71860
rect 1548 71851 1554 71854
rect 156 71814 162 71817
rect 126 71808 162 71814
rect 810 71814 816 71817
rect 810 71808 1584 71814
rect 126 71774 138 71808
rect 1572 71774 1584 71808
rect 126 71768 162 71774
rect 156 71765 162 71768
rect 810 71768 1584 71774
rect 810 71765 816 71768
rect 894 71728 900 71731
rect 126 71722 900 71728
rect 1548 71728 1554 71731
rect 1548 71722 1584 71728
rect 126 71688 138 71722
rect 1572 71688 1584 71722
rect 126 71682 900 71688
rect 894 71679 900 71682
rect 1548 71682 1584 71688
rect 1548 71679 1554 71682
rect 156 71642 162 71645
rect 126 71636 162 71642
rect 810 71642 816 71645
rect 810 71636 1584 71642
rect 126 71602 138 71636
rect 1572 71602 1584 71636
rect 126 71596 162 71602
rect 156 71593 162 71596
rect 810 71596 1584 71602
rect 810 71593 816 71596
rect 894 71556 900 71559
rect 126 71550 900 71556
rect 1548 71556 1554 71559
rect 1548 71550 1584 71556
rect 126 71516 138 71550
rect 1572 71516 1584 71550
rect 126 71510 900 71516
rect 894 71507 900 71510
rect 1548 71510 1584 71516
rect 1548 71507 1554 71510
rect 156 71470 162 71473
rect 126 71464 162 71470
rect 810 71470 816 71473
rect 810 71464 1584 71470
rect 126 71430 138 71464
rect 1572 71430 1584 71464
rect 126 71424 162 71430
rect 156 71421 162 71424
rect 810 71424 1584 71430
rect 810 71421 816 71424
rect 894 71384 900 71387
rect 126 71378 900 71384
rect 1548 71384 1554 71387
rect 1548 71378 1584 71384
rect 126 71344 138 71378
rect 1572 71344 1584 71378
rect 126 71338 900 71344
rect 894 71335 900 71338
rect 1548 71338 1584 71344
rect 1548 71335 1554 71338
rect 156 71298 162 71301
rect 126 71292 162 71298
rect 810 71298 816 71301
rect 810 71292 1584 71298
rect 126 71258 138 71292
rect 1572 71258 1584 71292
rect 126 71252 162 71258
rect 156 71249 162 71252
rect 810 71252 1584 71258
rect 810 71249 816 71252
rect 894 71212 900 71215
rect 126 71206 900 71212
rect 1548 71212 1554 71215
rect 1548 71206 1584 71212
rect 126 71172 138 71206
rect 1572 71172 1584 71206
rect 126 71166 900 71172
rect 894 71163 900 71166
rect 1548 71166 1584 71172
rect 1548 71163 1554 71166
rect 156 71126 162 71129
rect 126 71120 162 71126
rect 810 71126 816 71129
rect 810 71120 1584 71126
rect 126 71086 138 71120
rect 1572 71086 1584 71120
rect 126 71080 162 71086
rect 156 71077 162 71080
rect 810 71080 1584 71086
rect 810 71077 816 71080
rect 894 71040 900 71043
rect 126 71034 900 71040
rect 1548 71040 1554 71043
rect 1548 71034 1584 71040
rect 126 71000 138 71034
rect 1572 71000 1584 71034
rect 126 70994 900 71000
rect 894 70991 900 70994
rect 1548 70994 1584 71000
rect 1548 70991 1554 70994
rect 156 70954 162 70957
rect 126 70948 162 70954
rect 810 70954 816 70957
rect 810 70948 1584 70954
rect 126 70914 138 70948
rect 1572 70914 1584 70948
rect 126 70908 162 70914
rect 156 70905 162 70908
rect 810 70908 1584 70914
rect 810 70905 816 70908
rect 894 70868 900 70871
rect 126 70862 900 70868
rect 1548 70868 1554 70871
rect 1548 70862 1584 70868
rect 126 70828 138 70862
rect 1572 70828 1584 70862
rect 126 70822 900 70828
rect 894 70819 900 70822
rect 1548 70822 1584 70828
rect 1548 70819 1554 70822
rect 156 70782 162 70785
rect 126 70776 162 70782
rect 810 70782 816 70785
rect 810 70776 1584 70782
rect 126 70742 138 70776
rect 1572 70742 1584 70776
rect 126 70736 162 70742
rect 156 70733 162 70736
rect 810 70736 1584 70742
rect 810 70733 816 70736
rect 894 70696 900 70699
rect 126 70690 900 70696
rect 1548 70696 1554 70699
rect 1548 70690 1584 70696
rect 126 70656 138 70690
rect 1572 70656 1584 70690
rect 126 70650 900 70656
rect 894 70647 900 70650
rect 1548 70650 1584 70656
rect 1548 70647 1554 70650
rect 156 70610 162 70613
rect 126 70604 162 70610
rect 810 70610 816 70613
rect 810 70604 1584 70610
rect 126 70570 138 70604
rect 1572 70570 1584 70604
rect 126 70564 162 70570
rect 156 70561 162 70564
rect 810 70564 1584 70570
rect 810 70561 816 70564
rect 894 70524 900 70527
rect 126 70518 900 70524
rect 1548 70524 1554 70527
rect 1548 70518 1584 70524
rect 126 70484 138 70518
rect 1572 70484 1584 70518
rect 126 70478 900 70484
rect 894 70475 900 70478
rect 1548 70478 1584 70484
rect 1548 70475 1554 70478
rect 156 70438 162 70441
rect 126 70432 162 70438
rect 810 70438 816 70441
rect 810 70432 1584 70438
rect 126 70398 138 70432
rect 1572 70398 1584 70432
rect 126 70392 162 70398
rect 156 70389 162 70392
rect 810 70392 1584 70398
rect 810 70389 816 70392
rect 894 70352 900 70355
rect 126 70346 900 70352
rect 1548 70352 1554 70355
rect 1548 70346 1584 70352
rect 126 70312 138 70346
rect 1572 70312 1584 70346
rect 126 70306 900 70312
rect 894 70303 900 70306
rect 1548 70306 1584 70312
rect 1548 70303 1554 70306
rect 156 70266 162 70269
rect 126 70260 162 70266
rect 810 70266 816 70269
rect 810 70260 1584 70266
rect 126 70226 138 70260
rect 1572 70226 1584 70260
rect 126 70220 162 70226
rect 156 70217 162 70220
rect 810 70220 1584 70226
rect 810 70217 816 70220
rect 894 70180 900 70183
rect 126 70174 900 70180
rect 1548 70180 1554 70183
rect 1548 70174 1584 70180
rect 126 70140 138 70174
rect 1572 70140 1584 70174
rect 126 70134 900 70140
rect 894 70131 900 70134
rect 1548 70134 1584 70140
rect 1548 70131 1554 70134
rect 156 70094 162 70097
rect 126 70088 162 70094
rect 810 70094 816 70097
rect 810 70088 1584 70094
rect 126 70054 138 70088
rect 1572 70054 1584 70088
rect 126 70048 162 70054
rect 156 70045 162 70048
rect 810 70048 1584 70054
rect 810 70045 816 70048
rect 894 70008 900 70011
rect 126 70002 900 70008
rect 1548 70008 1554 70011
rect 1548 70002 1584 70008
rect 126 69968 138 70002
rect 1572 69968 1584 70002
rect 126 69962 900 69968
rect 894 69959 900 69962
rect 1548 69962 1584 69968
rect 1548 69959 1554 69962
rect 156 69922 162 69925
rect 126 69916 162 69922
rect 810 69922 816 69925
rect 810 69916 1584 69922
rect 126 69882 138 69916
rect 1572 69882 1584 69916
rect 126 69876 162 69882
rect 156 69873 162 69876
rect 810 69876 1584 69882
rect 810 69873 816 69876
rect 894 69836 900 69839
rect 126 69830 900 69836
rect 1548 69836 1554 69839
rect 1548 69830 1584 69836
rect 126 69796 138 69830
rect 1572 69796 1584 69830
rect 126 69790 900 69796
rect 894 69787 900 69790
rect 1548 69790 1584 69796
rect 1548 69787 1554 69790
rect 156 69750 162 69753
rect 126 69744 162 69750
rect 810 69750 816 69753
rect 810 69744 1584 69750
rect 126 69710 138 69744
rect 1572 69710 1584 69744
rect 126 69704 162 69710
rect 156 69701 162 69704
rect 810 69704 1584 69710
rect 810 69701 816 69704
rect 894 69664 900 69667
rect 126 69658 900 69664
rect 1548 69664 1554 69667
rect 1548 69658 1584 69664
rect 126 69624 138 69658
rect 1572 69624 1584 69658
rect 126 69618 900 69624
rect 894 69615 900 69618
rect 1548 69618 1584 69624
rect 1548 69615 1554 69618
rect 156 69578 162 69581
rect 126 69572 162 69578
rect 810 69578 816 69581
rect 810 69572 1584 69578
rect 126 69538 138 69572
rect 1572 69538 1584 69572
rect 126 69532 162 69538
rect 156 69529 162 69532
rect 810 69532 1584 69538
rect 810 69529 816 69532
rect 894 69492 900 69495
rect 126 69486 900 69492
rect 1548 69492 1554 69495
rect 1548 69486 1584 69492
rect 126 69452 138 69486
rect 1572 69452 1584 69486
rect 126 69446 900 69452
rect 894 69443 900 69446
rect 1548 69446 1584 69452
rect 1548 69443 1554 69446
rect 156 69406 162 69409
rect 126 69400 162 69406
rect 810 69406 816 69409
rect 810 69400 1584 69406
rect 126 69366 138 69400
rect 1572 69366 1584 69400
rect 126 69360 162 69366
rect 156 69357 162 69360
rect 810 69360 1584 69366
rect 810 69357 816 69360
rect 894 69320 900 69323
rect 126 69314 900 69320
rect 1548 69320 1554 69323
rect 1548 69314 1584 69320
rect 126 69280 138 69314
rect 1572 69280 1584 69314
rect 126 69274 900 69280
rect 894 69271 900 69274
rect 1548 69274 1584 69280
rect 1548 69271 1554 69274
rect 156 69234 162 69237
rect 126 69228 162 69234
rect 810 69234 816 69237
rect 810 69228 1584 69234
rect 126 69194 138 69228
rect 1572 69194 1584 69228
rect 126 69188 162 69194
rect 156 69185 162 69188
rect 810 69188 1584 69194
rect 810 69185 816 69188
rect 894 69148 900 69151
rect 126 69142 900 69148
rect 1548 69148 1554 69151
rect 1548 69142 1584 69148
rect 126 69108 138 69142
rect 1572 69108 1584 69142
rect 126 69102 900 69108
rect 894 69099 900 69102
rect 1548 69102 1584 69108
rect 1548 69099 1554 69102
rect 156 69062 162 69065
rect 126 69056 162 69062
rect 810 69062 816 69065
rect 810 69056 1584 69062
rect 126 69022 138 69056
rect 1572 69022 1584 69056
rect 126 69016 162 69022
rect 156 69013 162 69016
rect 810 69016 1584 69022
rect 810 69013 816 69016
rect 894 68976 900 68979
rect 126 68970 900 68976
rect 1548 68976 1554 68979
rect 1548 68970 1584 68976
rect 126 68936 138 68970
rect 1572 68936 1584 68970
rect 126 68930 900 68936
rect 894 68927 900 68930
rect 1548 68930 1584 68936
rect 1548 68927 1554 68930
rect 156 68890 162 68893
rect 126 68884 162 68890
rect 810 68890 816 68893
rect 810 68884 1584 68890
rect 126 68850 138 68884
rect 1572 68850 1584 68884
rect 126 68844 162 68850
rect 156 68841 162 68844
rect 810 68844 1584 68850
rect 810 68841 816 68844
rect 894 68804 900 68807
rect 126 68798 900 68804
rect 1548 68804 1554 68807
rect 1548 68798 1584 68804
rect 126 68764 138 68798
rect 1572 68764 1584 68798
rect 126 68758 900 68764
rect 894 68755 900 68758
rect 1548 68758 1584 68764
rect 1548 68755 1554 68758
rect 156 68718 162 68721
rect 126 68712 162 68718
rect 810 68718 816 68721
rect 810 68712 1584 68718
rect 126 68678 138 68712
rect 1572 68678 1584 68712
rect 126 68672 162 68678
rect 156 68669 162 68672
rect 810 68672 1584 68678
rect 810 68669 816 68672
rect 894 68632 900 68635
rect 126 68626 900 68632
rect 1548 68632 1554 68635
rect 1548 68626 1584 68632
rect 126 68592 138 68626
rect 1572 68592 1584 68626
rect 126 68586 900 68592
rect 894 68583 900 68586
rect 1548 68586 1584 68592
rect 1548 68583 1554 68586
rect 156 68546 162 68549
rect 126 68540 162 68546
rect 810 68546 816 68549
rect 810 68540 1584 68546
rect 126 68506 138 68540
rect 1572 68506 1584 68540
rect 126 68500 162 68506
rect 156 68497 162 68500
rect 810 68500 1584 68506
rect 810 68497 816 68500
rect 894 68460 900 68463
rect 126 68454 900 68460
rect 1548 68460 1554 68463
rect 1548 68454 1584 68460
rect 126 68420 138 68454
rect 1572 68420 1584 68454
rect 126 68414 900 68420
rect 894 68411 900 68414
rect 1548 68414 1584 68420
rect 1548 68411 1554 68414
rect 156 68374 162 68377
rect 126 68368 162 68374
rect 810 68374 816 68377
rect 810 68368 1584 68374
rect 126 68334 138 68368
rect 1572 68334 1584 68368
rect 126 68328 162 68334
rect 156 68325 162 68328
rect 810 68328 1584 68334
rect 810 68325 816 68328
rect 894 68288 900 68291
rect 126 68282 900 68288
rect 1548 68288 1554 68291
rect 1548 68282 1584 68288
rect 126 68248 138 68282
rect 1572 68248 1584 68282
rect 126 68242 900 68248
rect 894 68239 900 68242
rect 1548 68242 1584 68248
rect 1548 68239 1554 68242
rect 156 68202 162 68205
rect 126 68196 162 68202
rect 810 68202 816 68205
rect 810 68196 1584 68202
rect 126 68162 138 68196
rect 1572 68162 1584 68196
rect 126 68156 162 68162
rect 156 68153 162 68156
rect 810 68156 1584 68162
rect 810 68153 816 68156
rect 894 68116 900 68119
rect 126 68110 900 68116
rect 1548 68116 1554 68119
rect 1548 68110 1584 68116
rect 126 68076 138 68110
rect 1572 68076 1584 68110
rect 126 68070 900 68076
rect 894 68067 900 68070
rect 1548 68070 1584 68076
rect 1548 68067 1554 68070
rect 156 68030 162 68033
rect 126 68024 162 68030
rect 810 68030 816 68033
rect 810 68024 1584 68030
rect 126 67990 138 68024
rect 1572 67990 1584 68024
rect 126 67984 162 67990
rect 156 67981 162 67984
rect 810 67984 1584 67990
rect 810 67981 816 67984
rect 894 67944 900 67947
rect 126 67938 900 67944
rect 1548 67944 1554 67947
rect 1548 67938 1584 67944
rect 126 67904 138 67938
rect 1572 67904 1584 67938
rect 126 67898 900 67904
rect 894 67895 900 67898
rect 1548 67898 1584 67904
rect 1548 67895 1554 67898
rect 156 67858 162 67861
rect 126 67852 162 67858
rect 810 67858 816 67861
rect 810 67852 1584 67858
rect 126 67818 138 67852
rect 1572 67818 1584 67852
rect 126 67812 162 67818
rect 156 67809 162 67812
rect 810 67812 1584 67818
rect 810 67809 816 67812
rect 894 67772 900 67775
rect 126 67766 900 67772
rect 1548 67772 1554 67775
rect 1548 67766 1584 67772
rect 126 67732 138 67766
rect 1572 67732 1584 67766
rect 126 67726 900 67732
rect 894 67723 900 67726
rect 1548 67726 1584 67732
rect 1548 67723 1554 67726
rect 156 67686 162 67689
rect 126 67680 162 67686
rect 810 67686 816 67689
rect 810 67680 1584 67686
rect 126 67646 138 67680
rect 1572 67646 1584 67680
rect 126 67640 162 67646
rect 156 67637 162 67640
rect 810 67640 1584 67646
rect 810 67637 816 67640
rect 894 67600 900 67603
rect 126 67594 900 67600
rect 1548 67600 1554 67603
rect 1548 67594 1584 67600
rect 126 67560 138 67594
rect 1572 67560 1584 67594
rect 126 67554 900 67560
rect 894 67551 900 67554
rect 1548 67554 1584 67560
rect 1548 67551 1554 67554
rect 156 67514 162 67517
rect 126 67508 162 67514
rect 810 67514 816 67517
rect 810 67508 1584 67514
rect 126 67474 138 67508
rect 1572 67474 1584 67508
rect 126 67468 162 67474
rect 156 67465 162 67468
rect 810 67468 1584 67474
rect 810 67465 816 67468
rect 894 67428 900 67431
rect 126 67422 900 67428
rect 1548 67428 1554 67431
rect 1548 67422 1584 67428
rect 126 67388 138 67422
rect 1572 67388 1584 67422
rect 126 67382 900 67388
rect 894 67379 900 67382
rect 1548 67382 1584 67388
rect 1548 67379 1554 67382
rect 156 67342 162 67345
rect 126 67336 162 67342
rect 810 67342 816 67345
rect 810 67336 1584 67342
rect 126 67302 138 67336
rect 1572 67302 1584 67336
rect 126 67296 162 67302
rect 156 67293 162 67296
rect 810 67296 1584 67302
rect 810 67293 816 67296
rect 894 67256 900 67259
rect 126 67250 900 67256
rect 1548 67256 1554 67259
rect 1548 67250 1584 67256
rect 126 67216 138 67250
rect 1572 67216 1584 67250
rect 126 67210 900 67216
rect 894 67207 900 67210
rect 1548 67210 1584 67216
rect 1548 67207 1554 67210
rect 156 67170 162 67173
rect 126 67164 162 67170
rect 810 67170 816 67173
rect 810 67164 1584 67170
rect 126 67130 138 67164
rect 1572 67130 1584 67164
rect 126 67124 162 67130
rect 156 67121 162 67124
rect 810 67124 1584 67130
rect 810 67121 816 67124
rect 894 67084 900 67087
rect 126 67078 900 67084
rect 1548 67084 1554 67087
rect 1548 67078 1584 67084
rect 126 67044 138 67078
rect 1572 67044 1584 67078
rect 126 67038 900 67044
rect 894 67035 900 67038
rect 1548 67038 1584 67044
rect 1548 67035 1554 67038
rect 156 66998 162 67001
rect 126 66992 162 66998
rect 810 66998 816 67001
rect 810 66992 1584 66998
rect 126 66958 138 66992
rect 1572 66958 1584 66992
rect 126 66952 162 66958
rect 156 66949 162 66952
rect 810 66952 1584 66958
rect 810 66949 816 66952
rect 894 66912 900 66915
rect 126 66906 900 66912
rect 1548 66912 1554 66915
rect 1548 66906 1584 66912
rect 126 66872 138 66906
rect 1572 66872 1584 66906
rect 126 66866 900 66872
rect 894 66863 900 66866
rect 1548 66866 1584 66872
rect 1548 66863 1554 66866
rect 156 66826 162 66829
rect 126 66820 162 66826
rect 810 66826 816 66829
rect 810 66820 1584 66826
rect 126 66786 138 66820
rect 1572 66786 1584 66820
rect 126 66780 162 66786
rect 156 66777 162 66780
rect 810 66780 1584 66786
rect 810 66777 816 66780
rect 894 66740 900 66743
rect 126 66734 900 66740
rect 1548 66740 1554 66743
rect 1548 66734 1584 66740
rect 126 66700 138 66734
rect 1572 66700 1584 66734
rect 126 66694 900 66700
rect 894 66691 900 66694
rect 1548 66694 1584 66700
rect 1548 66691 1554 66694
rect 156 66654 162 66657
rect 126 66648 162 66654
rect 810 66654 816 66657
rect 810 66648 1584 66654
rect 126 66614 138 66648
rect 1572 66614 1584 66648
rect 126 66608 162 66614
rect 156 66605 162 66608
rect 810 66608 1584 66614
rect 810 66605 816 66608
rect 894 66568 900 66571
rect 126 66562 900 66568
rect 1548 66568 1554 66571
rect 1548 66562 1584 66568
rect 126 66528 138 66562
rect 1572 66528 1584 66562
rect 126 66522 900 66528
rect 894 66519 900 66522
rect 1548 66522 1584 66528
rect 1548 66519 1554 66522
rect 156 66482 162 66485
rect 126 66476 162 66482
rect 810 66482 816 66485
rect 810 66476 1584 66482
rect 126 66442 138 66476
rect 1572 66442 1584 66476
rect 126 66436 162 66442
rect 156 66433 162 66436
rect 810 66436 1584 66442
rect 810 66433 816 66436
rect 894 66396 900 66399
rect 126 66390 900 66396
rect 1548 66396 1554 66399
rect 1548 66390 1584 66396
rect 126 66356 138 66390
rect 1572 66356 1584 66390
rect 126 66350 900 66356
rect 894 66347 900 66350
rect 1548 66350 1584 66356
rect 1548 66347 1554 66350
rect 156 66310 162 66313
rect 126 66304 162 66310
rect 810 66310 816 66313
rect 810 66304 1584 66310
rect 126 66270 138 66304
rect 1572 66270 1584 66304
rect 126 66264 162 66270
rect 156 66261 162 66264
rect 810 66264 1584 66270
rect 810 66261 816 66264
rect 894 66224 900 66227
rect 126 66218 900 66224
rect 1548 66224 1554 66227
rect 1548 66218 1584 66224
rect 126 66184 138 66218
rect 1572 66184 1584 66218
rect 126 66178 900 66184
rect 894 66175 900 66178
rect 1548 66178 1584 66184
rect 1548 66175 1554 66178
rect 156 66138 162 66141
rect 126 66132 162 66138
rect 810 66138 816 66141
rect 810 66132 1584 66138
rect 126 66098 138 66132
rect 1572 66098 1584 66132
rect 126 66092 162 66098
rect 156 66089 162 66092
rect 810 66092 1584 66098
rect 810 66089 816 66092
rect 894 66052 900 66055
rect 126 66046 900 66052
rect 1548 66052 1554 66055
rect 1548 66046 1584 66052
rect 126 66012 138 66046
rect 1572 66012 1584 66046
rect 126 66006 900 66012
rect 894 66003 900 66006
rect 1548 66006 1584 66012
rect 1548 66003 1554 66006
rect 156 65966 162 65969
rect 126 65960 162 65966
rect 810 65966 816 65969
rect 810 65960 1584 65966
rect 126 65926 138 65960
rect 1572 65926 1584 65960
rect 126 65920 162 65926
rect 156 65917 162 65920
rect 810 65920 1584 65926
rect 810 65917 816 65920
rect 894 65880 900 65883
rect 126 65874 900 65880
rect 1548 65880 1554 65883
rect 1548 65874 1584 65880
rect 126 65840 138 65874
rect 1572 65840 1584 65874
rect 126 65834 900 65840
rect 894 65831 900 65834
rect 1548 65834 1584 65840
rect 1548 65831 1554 65834
rect 156 65794 162 65797
rect 126 65788 162 65794
rect 810 65794 816 65797
rect 810 65788 1584 65794
rect 126 65754 138 65788
rect 1572 65754 1584 65788
rect 126 65748 162 65754
rect 156 65745 162 65748
rect 810 65748 1584 65754
rect 810 65745 816 65748
rect 894 65708 900 65711
rect 126 65702 900 65708
rect 1548 65708 1554 65711
rect 1548 65702 1584 65708
rect 126 65668 138 65702
rect 1572 65668 1584 65702
rect 126 65662 900 65668
rect 894 65659 900 65662
rect 1548 65662 1584 65668
rect 1548 65659 1554 65662
rect 156 65622 162 65625
rect 126 65616 162 65622
rect 810 65622 816 65625
rect 810 65616 1584 65622
rect 126 65582 138 65616
rect 1572 65582 1584 65616
rect 126 65576 162 65582
rect 156 65573 162 65576
rect 810 65576 1584 65582
rect 810 65573 816 65576
rect 894 65536 900 65539
rect 126 65530 900 65536
rect 1548 65536 1554 65539
rect 1548 65530 1584 65536
rect 126 65496 138 65530
rect 1572 65496 1584 65530
rect 126 65490 900 65496
rect 894 65487 900 65490
rect 1548 65490 1584 65496
rect 1548 65487 1554 65490
rect 156 65450 162 65453
rect 126 65444 162 65450
rect 810 65450 816 65453
rect 810 65444 1584 65450
rect 126 65410 138 65444
rect 1572 65410 1584 65444
rect 126 65404 162 65410
rect 156 65401 162 65404
rect 810 65404 1584 65410
rect 810 65401 816 65404
rect 894 65364 900 65367
rect 126 65358 900 65364
rect 1548 65364 1554 65367
rect 1548 65358 1584 65364
rect 126 65324 138 65358
rect 1572 65324 1584 65358
rect 126 65318 900 65324
rect 894 65315 900 65318
rect 1548 65318 1584 65324
rect 1548 65315 1554 65318
rect 156 65278 162 65281
rect 126 65272 162 65278
rect 810 65278 816 65281
rect 810 65272 1584 65278
rect 126 65238 138 65272
rect 1572 65238 1584 65272
rect 126 65232 162 65238
rect 156 65229 162 65232
rect 810 65232 1584 65238
rect 810 65229 816 65232
rect 894 65192 900 65195
rect 126 65186 900 65192
rect 1548 65192 1554 65195
rect 1548 65186 1584 65192
rect 126 65152 138 65186
rect 1572 65152 1584 65186
rect 126 65146 900 65152
rect 894 65143 900 65146
rect 1548 65146 1584 65152
rect 1548 65143 1554 65146
rect 156 65106 162 65109
rect 126 65100 162 65106
rect 810 65106 816 65109
rect 810 65100 1584 65106
rect 126 65066 138 65100
rect 1572 65066 1584 65100
rect 126 65060 162 65066
rect 156 65057 162 65060
rect 810 65060 1584 65066
rect 810 65057 816 65060
rect 894 65020 900 65023
rect 126 65014 900 65020
rect 1548 65020 1554 65023
rect 1548 65014 1584 65020
rect 126 64980 138 65014
rect 1572 64980 1584 65014
rect 126 64974 900 64980
rect 894 64971 900 64974
rect 1548 64974 1584 64980
rect 1548 64971 1554 64974
rect 156 64934 162 64937
rect 126 64928 162 64934
rect 810 64934 816 64937
rect 810 64928 1584 64934
rect 126 64894 138 64928
rect 1572 64894 1584 64928
rect 126 64888 162 64894
rect 156 64885 162 64888
rect 810 64888 1584 64894
rect 810 64885 816 64888
rect 894 64848 900 64851
rect 126 64842 900 64848
rect 1548 64848 1554 64851
rect 1548 64842 1584 64848
rect 126 64808 138 64842
rect 1572 64808 1584 64842
rect 126 64802 900 64808
rect 894 64799 900 64802
rect 1548 64802 1584 64808
rect 1548 64799 1554 64802
rect 156 64762 162 64765
rect 126 64756 162 64762
rect 810 64762 816 64765
rect 810 64756 1584 64762
rect 126 64722 138 64756
rect 1572 64722 1584 64756
rect 126 64716 162 64722
rect 156 64713 162 64716
rect 810 64716 1584 64722
rect 810 64713 816 64716
rect 894 64676 900 64679
rect 126 64670 900 64676
rect 1548 64676 1554 64679
rect 1548 64670 1584 64676
rect 126 64636 138 64670
rect 1572 64636 1584 64670
rect 126 64630 900 64636
rect 894 64627 900 64630
rect 1548 64630 1584 64636
rect 1548 64627 1554 64630
rect 156 64590 162 64593
rect 126 64584 162 64590
rect 810 64590 816 64593
rect 810 64584 1584 64590
rect 126 64550 138 64584
rect 1572 64550 1584 64584
rect 126 64544 162 64550
rect 156 64541 162 64544
rect 810 64544 1584 64550
rect 810 64541 816 64544
rect 894 64504 900 64507
rect 126 64498 900 64504
rect 1548 64504 1554 64507
rect 1548 64498 1584 64504
rect 126 64464 138 64498
rect 1572 64464 1584 64498
rect 126 64458 900 64464
rect 894 64455 900 64458
rect 1548 64458 1584 64464
rect 1548 64455 1554 64458
rect 156 64418 162 64421
rect 126 64412 162 64418
rect 810 64418 816 64421
rect 810 64412 1584 64418
rect 126 64378 138 64412
rect 1572 64378 1584 64412
rect 126 64372 162 64378
rect 156 64369 162 64372
rect 810 64372 1584 64378
rect 810 64369 816 64372
rect 894 64332 900 64335
rect 126 64326 900 64332
rect 1548 64332 1554 64335
rect 1548 64326 1584 64332
rect 126 64292 138 64326
rect 1572 64292 1584 64326
rect 126 64286 900 64292
rect 894 64283 900 64286
rect 1548 64286 1584 64292
rect 1548 64283 1554 64286
rect 156 64246 162 64249
rect 126 64240 162 64246
rect 810 64246 816 64249
rect 810 64240 1584 64246
rect 126 64206 138 64240
rect 1572 64206 1584 64240
rect 126 64200 162 64206
rect 156 64197 162 64200
rect 810 64200 1584 64206
rect 810 64197 816 64200
rect 894 64160 900 64163
rect 126 64154 900 64160
rect 1548 64160 1554 64163
rect 1548 64154 1584 64160
rect 126 64120 138 64154
rect 1572 64120 1584 64154
rect 126 64114 900 64120
rect 894 64111 900 64114
rect 1548 64114 1584 64120
rect 1548 64111 1554 64114
rect 156 64074 162 64077
rect 126 64068 162 64074
rect 810 64074 816 64077
rect 810 64068 1584 64074
rect 126 64034 138 64068
rect 1572 64034 1584 64068
rect 126 64028 162 64034
rect 156 64025 162 64028
rect 810 64028 1584 64034
rect 810 64025 816 64028
rect 894 63988 900 63991
rect 126 63982 900 63988
rect 1548 63988 1554 63991
rect 1548 63982 1584 63988
rect 126 63948 138 63982
rect 1572 63948 1584 63982
rect 126 63942 900 63948
rect 894 63939 900 63942
rect 1548 63942 1584 63948
rect 1548 63939 1554 63942
rect 156 63902 162 63905
rect 126 63896 162 63902
rect 810 63902 816 63905
rect 810 63896 1584 63902
rect 126 63862 138 63896
rect 1572 63862 1584 63896
rect 126 63856 162 63862
rect 156 63853 162 63856
rect 810 63856 1584 63862
rect 810 63853 816 63856
rect 894 63816 900 63819
rect 126 63810 900 63816
rect 1548 63816 1554 63819
rect 1548 63810 1584 63816
rect 126 63776 138 63810
rect 1572 63776 1584 63810
rect 126 63770 900 63776
rect 894 63767 900 63770
rect 1548 63770 1584 63776
rect 1548 63767 1554 63770
rect 156 63730 162 63733
rect 126 63724 162 63730
rect 810 63730 816 63733
rect 810 63724 1584 63730
rect 126 63690 138 63724
rect 1572 63690 1584 63724
rect 126 63684 162 63690
rect 156 63681 162 63684
rect 810 63684 1584 63690
rect 810 63681 816 63684
rect 894 63644 900 63647
rect 126 63638 900 63644
rect 1548 63644 1554 63647
rect 1548 63638 1584 63644
rect 126 63604 138 63638
rect 1572 63604 1584 63638
rect 126 63598 900 63604
rect 894 63595 900 63598
rect 1548 63598 1584 63604
rect 1548 63595 1554 63598
rect 156 63558 162 63561
rect 126 63552 162 63558
rect 810 63558 816 63561
rect 810 63552 1584 63558
rect 126 63518 138 63552
rect 1572 63518 1584 63552
rect 126 63512 162 63518
rect 156 63509 162 63512
rect 810 63512 1584 63518
rect 810 63509 816 63512
rect 894 63472 900 63475
rect 126 63466 900 63472
rect 1548 63472 1554 63475
rect 1548 63466 1584 63472
rect 126 63432 138 63466
rect 1572 63432 1584 63466
rect 126 63426 900 63432
rect 894 63423 900 63426
rect 1548 63426 1584 63432
rect 1548 63423 1554 63426
rect 156 63386 162 63389
rect 126 63380 162 63386
rect 810 63386 816 63389
rect 810 63380 1584 63386
rect 126 63346 138 63380
rect 1572 63346 1584 63380
rect 126 63340 162 63346
rect 156 63337 162 63340
rect 810 63340 1584 63346
rect 810 63337 816 63340
rect 894 63300 900 63303
rect 126 63294 900 63300
rect 1548 63300 1554 63303
rect 1548 63294 1584 63300
rect 126 63260 138 63294
rect 1572 63260 1584 63294
rect 126 63254 900 63260
rect 894 63251 900 63254
rect 1548 63254 1584 63260
rect 1548 63251 1554 63254
rect 156 63214 162 63217
rect 126 63208 162 63214
rect 810 63214 816 63217
rect 810 63208 1584 63214
rect 126 63174 138 63208
rect 1572 63174 1584 63208
rect 126 63168 162 63174
rect 156 63165 162 63168
rect 810 63168 1584 63174
rect 810 63165 816 63168
rect 894 63128 900 63131
rect 126 63122 900 63128
rect 1548 63128 1554 63131
rect 1548 63122 1584 63128
rect 126 63088 138 63122
rect 1572 63088 1584 63122
rect 126 63082 900 63088
rect 894 63079 900 63082
rect 1548 63082 1584 63088
rect 1548 63079 1554 63082
rect 156 63042 162 63045
rect 126 63036 162 63042
rect 810 63042 816 63045
rect 810 63036 1584 63042
rect 126 63002 138 63036
rect 1572 63002 1584 63036
rect 126 62996 162 63002
rect 156 62993 162 62996
rect 810 62996 1584 63002
rect 810 62993 816 62996
rect 894 62956 900 62959
rect 126 62950 900 62956
rect 1548 62956 1554 62959
rect 1548 62950 1584 62956
rect 126 62916 138 62950
rect 1572 62916 1584 62950
rect 126 62910 900 62916
rect 894 62907 900 62910
rect 1548 62910 1584 62916
rect 1548 62907 1554 62910
rect 156 62870 162 62873
rect 126 62864 162 62870
rect 810 62870 816 62873
rect 810 62864 1584 62870
rect 126 62830 138 62864
rect 1572 62830 1584 62864
rect 126 62824 162 62830
rect 156 62821 162 62824
rect 810 62824 1584 62830
rect 810 62821 816 62824
rect 894 62784 900 62787
rect 126 62778 900 62784
rect 1548 62784 1554 62787
rect 1548 62778 1584 62784
rect 126 62744 138 62778
rect 1572 62744 1584 62778
rect 126 62738 900 62744
rect 894 62735 900 62738
rect 1548 62738 1584 62744
rect 1548 62735 1554 62738
rect 156 62698 162 62701
rect 126 62692 162 62698
rect 810 62698 816 62701
rect 810 62692 1584 62698
rect 126 62658 138 62692
rect 1572 62658 1584 62692
rect 126 62652 162 62658
rect 156 62649 162 62652
rect 810 62652 1584 62658
rect 810 62649 816 62652
rect 894 62612 900 62615
rect 126 62606 900 62612
rect 1548 62612 1554 62615
rect 1548 62606 1584 62612
rect 126 62572 138 62606
rect 1572 62572 1584 62606
rect 126 62566 900 62572
rect 894 62563 900 62566
rect 1548 62566 1584 62572
rect 1548 62563 1554 62566
rect 156 62526 162 62529
rect 126 62520 162 62526
rect 810 62526 816 62529
rect 810 62520 1584 62526
rect 126 62486 138 62520
rect 1572 62486 1584 62520
rect 126 62480 162 62486
rect 156 62477 162 62480
rect 810 62480 1584 62486
rect 810 62477 816 62480
rect 894 62440 900 62443
rect 126 62434 900 62440
rect 1548 62440 1554 62443
rect 1548 62434 1584 62440
rect 126 62400 138 62434
rect 1572 62400 1584 62434
rect 126 62394 900 62400
rect 894 62391 900 62394
rect 1548 62394 1584 62400
rect 1548 62391 1554 62394
rect 156 62354 162 62357
rect 126 62348 162 62354
rect 810 62354 816 62357
rect 810 62348 1584 62354
rect 126 62314 138 62348
rect 1572 62314 1584 62348
rect 126 62308 162 62314
rect 156 62305 162 62308
rect 810 62308 1584 62314
rect 810 62305 816 62308
rect 894 62268 900 62271
rect 126 62262 900 62268
rect 1548 62268 1554 62271
rect 1548 62262 1584 62268
rect 126 62228 138 62262
rect 1572 62228 1584 62262
rect 126 62222 900 62228
rect 894 62219 900 62222
rect 1548 62222 1584 62228
rect 1548 62219 1554 62222
rect 156 62182 162 62185
rect 126 62176 162 62182
rect 810 62182 816 62185
rect 810 62176 1584 62182
rect 126 62142 138 62176
rect 1572 62142 1584 62176
rect 126 62136 162 62142
rect 156 62133 162 62136
rect 810 62136 1584 62142
rect 810 62133 816 62136
rect 894 62096 900 62099
rect 126 62090 900 62096
rect 1548 62096 1554 62099
rect 1548 62090 1584 62096
rect 126 62056 138 62090
rect 1572 62056 1584 62090
rect 126 62050 900 62056
rect 894 62047 900 62050
rect 1548 62050 1584 62056
rect 1548 62047 1554 62050
rect 156 62010 162 62013
rect 126 62004 162 62010
rect 810 62010 816 62013
rect 810 62004 1584 62010
rect 126 61970 138 62004
rect 1572 61970 1584 62004
rect 126 61964 162 61970
rect 156 61961 162 61964
rect 810 61964 1584 61970
rect 810 61961 816 61964
rect 894 61924 900 61927
rect 126 61918 900 61924
rect 1548 61924 1554 61927
rect 1548 61918 1584 61924
rect 126 61884 138 61918
rect 1572 61884 1584 61918
rect 126 61878 900 61884
rect 894 61875 900 61878
rect 1548 61878 1584 61884
rect 1548 61875 1554 61878
rect 156 61838 162 61841
rect 126 61832 162 61838
rect 810 61838 816 61841
rect 810 61832 1584 61838
rect 126 61798 138 61832
rect 1572 61798 1584 61832
rect 126 61792 162 61798
rect 156 61789 162 61792
rect 810 61792 1584 61798
rect 810 61789 816 61792
rect 894 61752 900 61755
rect 126 61746 900 61752
rect 1548 61752 1554 61755
rect 1548 61746 1584 61752
rect 126 61712 138 61746
rect 1572 61712 1584 61746
rect 126 61706 900 61712
rect 894 61703 900 61706
rect 1548 61706 1584 61712
rect 1548 61703 1554 61706
rect 156 61666 162 61669
rect 126 61660 162 61666
rect 810 61666 816 61669
rect 810 61660 1584 61666
rect 126 61626 138 61660
rect 1572 61626 1584 61660
rect 126 61620 162 61626
rect 156 61617 162 61620
rect 810 61620 1584 61626
rect 810 61617 816 61620
rect 894 61580 900 61583
rect 126 61574 900 61580
rect 1548 61580 1554 61583
rect 1548 61574 1584 61580
rect 126 61540 138 61574
rect 1572 61540 1584 61574
rect 126 61534 900 61540
rect 894 61531 900 61534
rect 1548 61534 1584 61540
rect 1548 61531 1554 61534
rect 156 61494 162 61497
rect 126 61488 162 61494
rect 810 61494 816 61497
rect 810 61488 1584 61494
rect 126 61454 138 61488
rect 1572 61454 1584 61488
rect 126 61448 162 61454
rect 156 61445 162 61448
rect 810 61448 1584 61454
rect 810 61445 816 61448
rect 894 61408 900 61411
rect 126 61402 900 61408
rect 1548 61408 1554 61411
rect 1548 61402 1584 61408
rect 126 61368 138 61402
rect 1572 61368 1584 61402
rect 126 61362 900 61368
rect 894 61359 900 61362
rect 1548 61362 1584 61368
rect 1548 61359 1554 61362
rect 156 61322 162 61325
rect 126 61316 162 61322
rect 810 61322 816 61325
rect 810 61316 1584 61322
rect 126 61282 138 61316
rect 1572 61282 1584 61316
rect 126 61276 162 61282
rect 156 61273 162 61276
rect 810 61276 1584 61282
rect 810 61273 816 61276
rect 894 61236 900 61239
rect 126 61230 900 61236
rect 1548 61236 1554 61239
rect 1548 61230 1584 61236
rect 126 61196 138 61230
rect 1572 61196 1584 61230
rect 126 61190 900 61196
rect 894 61187 900 61190
rect 1548 61190 1584 61196
rect 1548 61187 1554 61190
rect 156 61150 162 61153
rect 126 61144 162 61150
rect 810 61150 816 61153
rect 810 61144 1584 61150
rect 126 61110 138 61144
rect 1572 61110 1584 61144
rect 126 61104 162 61110
rect 156 61101 162 61104
rect 810 61104 1584 61110
rect 810 61101 816 61104
rect 894 61064 900 61067
rect 126 61058 900 61064
rect 1548 61064 1554 61067
rect 1548 61058 1584 61064
rect 126 61024 138 61058
rect 1572 61024 1584 61058
rect 126 61018 900 61024
rect 894 61015 900 61018
rect 1548 61018 1584 61024
rect 1548 61015 1554 61018
rect 156 60978 162 60981
rect 126 60972 162 60978
rect 810 60978 816 60981
rect 810 60972 1584 60978
rect 126 60938 138 60972
rect 1572 60938 1584 60972
rect 126 60932 162 60938
rect 156 60929 162 60932
rect 810 60932 1584 60938
rect 810 60929 816 60932
rect 894 60892 900 60895
rect 126 60886 900 60892
rect 1548 60892 1554 60895
rect 1548 60886 1584 60892
rect 126 60852 138 60886
rect 1572 60852 1584 60886
rect 126 60846 900 60852
rect 894 60843 900 60846
rect 1548 60846 1584 60852
rect 1548 60843 1554 60846
rect 156 60806 162 60809
rect 126 60800 162 60806
rect 810 60806 816 60809
rect 810 60800 1584 60806
rect 126 60766 138 60800
rect 1572 60766 1584 60800
rect 126 60760 162 60766
rect 156 60757 162 60760
rect 810 60760 1584 60766
rect 810 60757 816 60760
rect 894 60720 900 60723
rect 126 60714 900 60720
rect 1548 60720 1554 60723
rect 1548 60714 1584 60720
rect 126 60680 138 60714
rect 1572 60680 1584 60714
rect 126 60674 900 60680
rect 894 60671 900 60674
rect 1548 60674 1584 60680
rect 1548 60671 1554 60674
rect 156 60634 162 60637
rect 126 60628 162 60634
rect 810 60634 816 60637
rect 810 60628 1584 60634
rect 126 60594 138 60628
rect 1572 60594 1584 60628
rect 126 60588 162 60594
rect 156 60585 162 60588
rect 810 60588 1584 60594
rect 810 60585 816 60588
rect 894 60548 900 60551
rect 126 60542 900 60548
rect 1548 60548 1554 60551
rect 1548 60542 1584 60548
rect 126 60508 138 60542
rect 1572 60508 1584 60542
rect 126 60502 900 60508
rect 894 60499 900 60502
rect 1548 60502 1584 60508
rect 1548 60499 1554 60502
rect 156 60462 162 60465
rect 126 60456 162 60462
rect 810 60462 816 60465
rect 810 60456 1584 60462
rect 126 60422 138 60456
rect 1572 60422 1584 60456
rect 126 60416 162 60422
rect 156 60413 162 60416
rect 810 60416 1584 60422
rect 810 60413 816 60416
rect 894 60376 900 60379
rect 126 60370 900 60376
rect 1548 60376 1554 60379
rect 1548 60370 1584 60376
rect 126 60336 138 60370
rect 1572 60336 1584 60370
rect 126 60330 900 60336
rect 894 60327 900 60330
rect 1548 60330 1584 60336
rect 1548 60327 1554 60330
rect 156 60290 162 60293
rect 126 60284 162 60290
rect 810 60290 816 60293
rect 810 60284 1584 60290
rect 126 60250 138 60284
rect 1572 60250 1584 60284
rect 126 60244 162 60250
rect 156 60241 162 60244
rect 810 60244 1584 60250
rect 810 60241 816 60244
rect 894 60204 900 60207
rect 126 60198 900 60204
rect 1548 60204 1554 60207
rect 1548 60198 1584 60204
rect 126 60164 138 60198
rect 1572 60164 1584 60198
rect 126 60158 900 60164
rect 894 60155 900 60158
rect 1548 60158 1584 60164
rect 1548 60155 1554 60158
rect 156 60118 162 60121
rect 126 60112 162 60118
rect 810 60118 816 60121
rect 810 60112 1584 60118
rect 126 60078 138 60112
rect 1572 60078 1584 60112
rect 126 60072 162 60078
rect 156 60069 162 60072
rect 810 60072 1584 60078
rect 810 60069 816 60072
rect 894 60032 900 60035
rect 126 60026 900 60032
rect 1548 60032 1554 60035
rect 1548 60026 1584 60032
rect 126 59992 138 60026
rect 1572 59992 1584 60026
rect 126 59986 900 59992
rect 894 59983 900 59986
rect 1548 59986 1584 59992
rect 1548 59983 1554 59986
rect 156 59946 162 59949
rect 126 59940 162 59946
rect 810 59946 816 59949
rect 810 59940 1584 59946
rect 126 59906 138 59940
rect 1572 59906 1584 59940
rect 126 59900 162 59906
rect 156 59897 162 59900
rect 810 59900 1584 59906
rect 810 59897 816 59900
rect 894 59860 900 59863
rect 126 59854 900 59860
rect 1548 59860 1554 59863
rect 1548 59854 1584 59860
rect 126 59820 138 59854
rect 1572 59820 1584 59854
rect 126 59814 900 59820
rect 894 59811 900 59814
rect 1548 59814 1584 59820
rect 1548 59811 1554 59814
rect 156 59774 162 59777
rect 126 59768 162 59774
rect 810 59774 816 59777
rect 810 59768 1584 59774
rect 126 59734 138 59768
rect 1572 59734 1584 59768
rect 126 59728 162 59734
rect 156 59725 162 59728
rect 810 59728 1584 59734
rect 810 59725 816 59728
rect 894 59688 900 59691
rect 126 59682 900 59688
rect 1548 59688 1554 59691
rect 1548 59682 1584 59688
rect 126 59648 138 59682
rect 1572 59648 1584 59682
rect 126 59642 900 59648
rect 894 59639 900 59642
rect 1548 59642 1584 59648
rect 1548 59639 1554 59642
rect 156 59602 162 59605
rect 126 59596 162 59602
rect 810 59602 816 59605
rect 810 59596 1584 59602
rect 126 59562 138 59596
rect 1572 59562 1584 59596
rect 126 59556 162 59562
rect 156 59553 162 59556
rect 810 59556 1584 59562
rect 810 59553 816 59556
rect 894 59516 900 59519
rect 126 59510 900 59516
rect 1548 59516 1554 59519
rect 1548 59510 1584 59516
rect 126 59476 138 59510
rect 1572 59476 1584 59510
rect 126 59470 900 59476
rect 894 59467 900 59470
rect 1548 59470 1584 59476
rect 1548 59467 1554 59470
rect 156 59430 162 59433
rect 126 59424 162 59430
rect 810 59430 816 59433
rect 810 59424 1584 59430
rect 126 59390 138 59424
rect 1572 59390 1584 59424
rect 126 59384 162 59390
rect 156 59381 162 59384
rect 810 59384 1584 59390
rect 810 59381 816 59384
rect 894 59344 900 59347
rect 126 59338 900 59344
rect 1548 59344 1554 59347
rect 1548 59338 1584 59344
rect 126 59304 138 59338
rect 1572 59304 1584 59338
rect 126 59298 900 59304
rect 894 59295 900 59298
rect 1548 59298 1584 59304
rect 1548 59295 1554 59298
rect 156 59258 162 59261
rect 126 59252 162 59258
rect 810 59258 816 59261
rect 810 59252 1584 59258
rect 126 59218 138 59252
rect 1572 59218 1584 59252
rect 126 59212 162 59218
rect 156 59209 162 59212
rect 810 59212 1584 59218
rect 810 59209 816 59212
rect 894 59172 900 59175
rect 126 59166 900 59172
rect 1548 59172 1554 59175
rect 1548 59166 1584 59172
rect 126 59132 138 59166
rect 1572 59132 1584 59166
rect 126 59126 900 59132
rect 894 59123 900 59126
rect 1548 59126 1584 59132
rect 1548 59123 1554 59126
rect 156 59086 162 59089
rect 126 59080 162 59086
rect 810 59086 816 59089
rect 810 59080 1584 59086
rect 126 59046 138 59080
rect 1572 59046 1584 59080
rect 126 59040 162 59046
rect 156 59037 162 59040
rect 810 59040 1584 59046
rect 810 59037 816 59040
rect 894 59000 900 59003
rect 126 58994 900 59000
rect 1548 59000 1554 59003
rect 1548 58994 1584 59000
rect 126 58960 138 58994
rect 1572 58960 1584 58994
rect 126 58954 900 58960
rect 894 58951 900 58954
rect 1548 58954 1584 58960
rect 1548 58951 1554 58954
rect 156 58914 162 58917
rect 126 58908 162 58914
rect 810 58914 816 58917
rect 810 58908 1584 58914
rect 126 58874 138 58908
rect 1572 58874 1584 58908
rect 126 58868 162 58874
rect 156 58865 162 58868
rect 810 58868 1584 58874
rect 810 58865 816 58868
rect 894 58828 900 58831
rect 126 58822 900 58828
rect 1548 58828 1554 58831
rect 1548 58822 1584 58828
rect 126 58788 138 58822
rect 1572 58788 1584 58822
rect 126 58782 900 58788
rect 894 58779 900 58782
rect 1548 58782 1584 58788
rect 1548 58779 1554 58782
rect 156 58742 162 58745
rect 126 58736 162 58742
rect 810 58742 816 58745
rect 810 58736 1584 58742
rect 126 58702 138 58736
rect 1572 58702 1584 58736
rect 126 58696 162 58702
rect 156 58693 162 58696
rect 810 58696 1584 58702
rect 810 58693 816 58696
rect 894 58656 900 58659
rect 126 58650 900 58656
rect 1548 58656 1554 58659
rect 1548 58650 1584 58656
rect 126 58616 138 58650
rect 1572 58616 1584 58650
rect 126 58610 900 58616
rect 894 58607 900 58610
rect 1548 58610 1584 58616
rect 1548 58607 1554 58610
rect 156 58570 162 58573
rect 126 58564 162 58570
rect 810 58570 816 58573
rect 810 58564 1584 58570
rect 126 58530 138 58564
rect 1572 58530 1584 58564
rect 126 58524 162 58530
rect 156 58521 162 58524
rect 810 58524 1584 58530
rect 810 58521 816 58524
rect 894 58484 900 58487
rect 126 58478 900 58484
rect 1548 58484 1554 58487
rect 1548 58478 1584 58484
rect 126 58444 138 58478
rect 1572 58444 1584 58478
rect 126 58438 900 58444
rect 894 58435 900 58438
rect 1548 58438 1584 58444
rect 1548 58435 1554 58438
rect 156 58398 162 58401
rect 126 58392 162 58398
rect 810 58398 816 58401
rect 810 58392 1584 58398
rect 126 58358 138 58392
rect 1572 58358 1584 58392
rect 126 58352 162 58358
rect 156 58349 162 58352
rect 810 58352 1584 58358
rect 810 58349 816 58352
rect 894 58312 900 58315
rect 126 58306 900 58312
rect 1548 58312 1554 58315
rect 1548 58306 1584 58312
rect 126 58272 138 58306
rect 1572 58272 1584 58306
rect 126 58266 900 58272
rect 894 58263 900 58266
rect 1548 58266 1584 58272
rect 1548 58263 1554 58266
rect 156 58226 162 58229
rect 126 58220 162 58226
rect 810 58226 816 58229
rect 810 58220 1584 58226
rect 126 58186 138 58220
rect 1572 58186 1584 58220
rect 126 58180 162 58186
rect 156 58177 162 58180
rect 810 58180 1584 58186
rect 810 58177 816 58180
rect 894 58140 900 58143
rect 126 58134 900 58140
rect 1548 58140 1554 58143
rect 1548 58134 1584 58140
rect 126 58100 138 58134
rect 1572 58100 1584 58134
rect 126 58094 900 58100
rect 894 58091 900 58094
rect 1548 58094 1584 58100
rect 1548 58091 1554 58094
rect 156 58054 162 58057
rect 126 58048 162 58054
rect 810 58054 816 58057
rect 810 58048 1584 58054
rect 126 58014 138 58048
rect 1572 58014 1584 58048
rect 126 58008 162 58014
rect 156 58005 162 58008
rect 810 58008 1584 58014
rect 810 58005 816 58008
rect 894 57968 900 57971
rect 126 57962 900 57968
rect 1548 57968 1554 57971
rect 1548 57962 1584 57968
rect 126 57928 138 57962
rect 1572 57928 1584 57962
rect 126 57922 900 57928
rect 894 57919 900 57922
rect 1548 57922 1584 57928
rect 1548 57919 1554 57922
rect 156 57882 162 57885
rect 126 57876 162 57882
rect 810 57882 816 57885
rect 810 57876 1584 57882
rect 126 57842 138 57876
rect 1572 57842 1584 57876
rect 126 57836 162 57842
rect 156 57833 162 57836
rect 810 57836 1584 57842
rect 810 57833 816 57836
rect 894 57796 900 57799
rect 126 57790 900 57796
rect 1548 57796 1554 57799
rect 1548 57790 1584 57796
rect 126 57756 138 57790
rect 1572 57756 1584 57790
rect 126 57750 900 57756
rect 894 57747 900 57750
rect 1548 57750 1584 57756
rect 1548 57747 1554 57750
rect 156 57710 162 57713
rect 126 57704 162 57710
rect 810 57710 816 57713
rect 810 57704 1584 57710
rect 126 57670 138 57704
rect 1572 57670 1584 57704
rect 126 57664 162 57670
rect 156 57661 162 57664
rect 810 57664 1584 57670
rect 810 57661 816 57664
rect 894 57624 900 57627
rect 126 57618 900 57624
rect 1548 57624 1554 57627
rect 1548 57618 1584 57624
rect 126 57584 138 57618
rect 1572 57584 1584 57618
rect 126 57578 900 57584
rect 894 57575 900 57578
rect 1548 57578 1584 57584
rect 1548 57575 1554 57578
rect 156 57538 162 57541
rect 126 57532 162 57538
rect 810 57538 816 57541
rect 810 57532 1584 57538
rect 126 57498 138 57532
rect 1572 57498 1584 57532
rect 126 57492 162 57498
rect 156 57489 162 57492
rect 810 57492 1584 57498
rect 810 57489 816 57492
rect 894 57452 900 57455
rect 126 57446 900 57452
rect 1548 57452 1554 57455
rect 1548 57446 1584 57452
rect 126 57412 138 57446
rect 1572 57412 1584 57446
rect 126 57406 900 57412
rect 894 57403 900 57406
rect 1548 57406 1584 57412
rect 1548 57403 1554 57406
rect 156 57366 162 57369
rect 126 57360 162 57366
rect 810 57366 816 57369
rect 810 57360 1584 57366
rect 126 57326 138 57360
rect 1572 57326 1584 57360
rect 126 57320 162 57326
rect 156 57317 162 57320
rect 810 57320 1584 57326
rect 810 57317 816 57320
rect 894 57280 900 57283
rect 126 57274 900 57280
rect 1548 57280 1554 57283
rect 1548 57274 1584 57280
rect 126 57240 138 57274
rect 1572 57240 1584 57274
rect 126 57234 900 57240
rect 894 57231 900 57234
rect 1548 57234 1584 57240
rect 1548 57231 1554 57234
rect 156 57194 162 57197
rect 126 57188 162 57194
rect 810 57194 816 57197
rect 810 57188 1584 57194
rect 126 57154 138 57188
rect 1572 57154 1584 57188
rect 126 57148 162 57154
rect 156 57145 162 57148
rect 810 57148 1584 57154
rect 810 57145 816 57148
rect 894 57108 900 57111
rect 126 57102 900 57108
rect 1548 57108 1554 57111
rect 1548 57102 1584 57108
rect 126 57068 138 57102
rect 1572 57068 1584 57102
rect 126 57062 900 57068
rect 894 57059 900 57062
rect 1548 57062 1584 57068
rect 1548 57059 1554 57062
rect 156 57022 162 57025
rect 126 57016 162 57022
rect 810 57022 816 57025
rect 810 57016 1584 57022
rect 126 56982 138 57016
rect 1572 56982 1584 57016
rect 126 56976 162 56982
rect 156 56973 162 56976
rect 810 56976 1584 56982
rect 810 56973 816 56976
rect 894 56936 900 56939
rect 126 56930 900 56936
rect 1548 56936 1554 56939
rect 1548 56930 1584 56936
rect 126 56896 138 56930
rect 1572 56896 1584 56930
rect 126 56890 900 56896
rect 894 56887 900 56890
rect 1548 56890 1584 56896
rect 1548 56887 1554 56890
rect 156 56850 162 56853
rect 126 56844 162 56850
rect 810 56850 816 56853
rect 810 56844 1584 56850
rect 126 56810 138 56844
rect 1572 56810 1584 56844
rect 126 56804 162 56810
rect 156 56801 162 56804
rect 810 56804 1584 56810
rect 810 56801 816 56804
rect 894 56764 900 56767
rect 126 56758 900 56764
rect 1548 56764 1554 56767
rect 1548 56758 1584 56764
rect 126 56724 138 56758
rect 1572 56724 1584 56758
rect 126 56718 900 56724
rect 894 56715 900 56718
rect 1548 56718 1584 56724
rect 1548 56715 1554 56718
rect 156 56678 162 56681
rect 126 56672 162 56678
rect 810 56678 816 56681
rect 810 56672 1584 56678
rect 126 56638 138 56672
rect 1572 56638 1584 56672
rect 126 56632 162 56638
rect 156 56629 162 56632
rect 810 56632 1584 56638
rect 810 56629 816 56632
rect 894 56592 900 56595
rect 126 56586 900 56592
rect 1548 56592 1554 56595
rect 1548 56586 1584 56592
rect 126 56552 138 56586
rect 1572 56552 1584 56586
rect 126 56546 900 56552
rect 894 56543 900 56546
rect 1548 56546 1584 56552
rect 1548 56543 1554 56546
rect 156 56506 162 56509
rect 126 56500 162 56506
rect 810 56506 816 56509
rect 810 56500 1584 56506
rect 126 56466 138 56500
rect 1572 56466 1584 56500
rect 126 56460 162 56466
rect 156 56457 162 56460
rect 810 56460 1584 56466
rect 810 56457 816 56460
rect 894 56420 900 56423
rect 126 56414 900 56420
rect 1548 56420 1554 56423
rect 1548 56414 1584 56420
rect 126 56380 138 56414
rect 1572 56380 1584 56414
rect 126 56374 900 56380
rect 894 56371 900 56374
rect 1548 56374 1584 56380
rect 1548 56371 1554 56374
rect 156 56334 162 56337
rect 126 56328 162 56334
rect 810 56334 816 56337
rect 810 56328 1584 56334
rect 126 56294 138 56328
rect 1572 56294 1584 56328
rect 126 56288 162 56294
rect 156 56285 162 56288
rect 810 56288 1584 56294
rect 810 56285 816 56288
rect 894 56248 900 56251
rect 126 56242 900 56248
rect 1548 56248 1554 56251
rect 1548 56242 1584 56248
rect 126 56208 138 56242
rect 1572 56208 1584 56242
rect 126 56202 900 56208
rect 894 56199 900 56202
rect 1548 56202 1584 56208
rect 1548 56199 1554 56202
rect 156 56162 162 56165
rect 126 56156 162 56162
rect 810 56162 816 56165
rect 810 56156 1584 56162
rect 126 56122 138 56156
rect 1572 56122 1584 56156
rect 126 56116 162 56122
rect 156 56113 162 56116
rect 810 56116 1584 56122
rect 810 56113 816 56116
rect 894 56076 900 56079
rect 126 56070 900 56076
rect 1548 56076 1554 56079
rect 1548 56070 1584 56076
rect 126 56036 138 56070
rect 1572 56036 1584 56070
rect 126 56030 900 56036
rect 894 56027 900 56030
rect 1548 56030 1584 56036
rect 1548 56027 1554 56030
rect 156 55990 162 55993
rect 126 55984 162 55990
rect 810 55990 816 55993
rect 810 55984 1584 55990
rect 126 55950 138 55984
rect 1572 55950 1584 55984
rect 126 55944 162 55950
rect 156 55941 162 55944
rect 810 55944 1584 55950
rect 810 55941 816 55944
rect 894 55904 900 55907
rect 126 55898 900 55904
rect 1548 55904 1554 55907
rect 1548 55898 1584 55904
rect 126 55864 138 55898
rect 1572 55864 1584 55898
rect 126 55858 900 55864
rect 894 55855 900 55858
rect 1548 55858 1584 55864
rect 1548 55855 1554 55858
rect 156 55818 162 55821
rect 126 55812 162 55818
rect 810 55818 816 55821
rect 810 55812 1584 55818
rect 126 55778 138 55812
rect 1572 55778 1584 55812
rect 126 55772 162 55778
rect 156 55769 162 55772
rect 810 55772 1584 55778
rect 810 55769 816 55772
rect 894 55732 900 55735
rect 126 55726 900 55732
rect 1548 55732 1554 55735
rect 1548 55726 1584 55732
rect 126 55692 138 55726
rect 1572 55692 1584 55726
rect 126 55686 900 55692
rect 894 55683 900 55686
rect 1548 55686 1584 55692
rect 1548 55683 1554 55686
rect 156 55646 162 55649
rect 126 55640 162 55646
rect 810 55646 816 55649
rect 810 55640 1584 55646
rect 126 55606 138 55640
rect 1572 55606 1584 55640
rect 126 55600 162 55606
rect 156 55597 162 55600
rect 810 55600 1584 55606
rect 810 55597 816 55600
rect 894 55560 900 55563
rect 126 55554 900 55560
rect 1548 55560 1554 55563
rect 1548 55554 1584 55560
rect 126 55520 138 55554
rect 1572 55520 1584 55554
rect 126 55514 900 55520
rect 894 55511 900 55514
rect 1548 55514 1584 55520
rect 1548 55511 1554 55514
rect 156 55474 162 55477
rect 126 55468 162 55474
rect 810 55474 816 55477
rect 810 55468 1584 55474
rect 126 55434 138 55468
rect 1572 55434 1584 55468
rect 126 55428 162 55434
rect 156 55425 162 55428
rect 810 55428 1584 55434
rect 810 55425 816 55428
rect 894 55388 900 55391
rect 126 55382 900 55388
rect 1548 55388 1554 55391
rect 1548 55382 1584 55388
rect 126 55348 138 55382
rect 1572 55348 1584 55382
rect 126 55342 900 55348
rect 894 55339 900 55342
rect 1548 55342 1584 55348
rect 1548 55339 1554 55342
rect 156 55302 162 55305
rect 126 55296 162 55302
rect 810 55302 816 55305
rect 810 55296 1584 55302
rect 126 55262 138 55296
rect 1572 55262 1584 55296
rect 126 55256 162 55262
rect 156 55253 162 55256
rect 810 55256 1584 55262
rect 810 55253 816 55256
rect 894 55216 900 55219
rect 126 55210 900 55216
rect 1548 55216 1554 55219
rect 1548 55210 1584 55216
rect 126 55176 138 55210
rect 1572 55176 1584 55210
rect 126 55170 900 55176
rect 894 55167 900 55170
rect 1548 55170 1584 55176
rect 1548 55167 1554 55170
rect 156 55130 162 55133
rect 126 55124 162 55130
rect 810 55130 816 55133
rect 810 55124 1584 55130
rect 126 55090 138 55124
rect 1572 55090 1584 55124
rect 126 55084 162 55090
rect 156 55081 162 55084
rect 810 55084 1584 55090
rect 810 55081 816 55084
rect 894 55044 900 55047
rect 126 55038 900 55044
rect 1548 55044 1554 55047
rect 1548 55038 1584 55044
rect 126 55004 138 55038
rect 1572 55004 1584 55038
rect 126 54998 900 55004
rect 894 54995 900 54998
rect 1548 54998 1584 55004
rect 1548 54995 1554 54998
rect 156 54958 162 54961
rect 126 54952 162 54958
rect 810 54958 816 54961
rect 810 54952 1584 54958
rect 126 54918 138 54952
rect 1572 54918 1584 54952
rect 126 54912 162 54918
rect 156 54909 162 54912
rect 810 54912 1584 54918
rect 810 54909 816 54912
rect 894 54872 900 54875
rect 126 54866 900 54872
rect 1548 54872 1554 54875
rect 1548 54866 1584 54872
rect 126 54832 138 54866
rect 1572 54832 1584 54866
rect 126 54826 900 54832
rect 894 54823 900 54826
rect 1548 54826 1584 54832
rect 1548 54823 1554 54826
rect 156 54786 162 54789
rect 126 54780 162 54786
rect 810 54786 816 54789
rect 810 54780 1584 54786
rect 126 54746 138 54780
rect 1572 54746 1584 54780
rect 126 54740 162 54746
rect 156 54737 162 54740
rect 810 54740 1584 54746
rect 810 54737 816 54740
rect 894 54700 900 54703
rect 126 54694 900 54700
rect 1548 54700 1554 54703
rect 1548 54694 1584 54700
rect 126 54660 138 54694
rect 1572 54660 1584 54694
rect 126 54654 900 54660
rect 894 54651 900 54654
rect 1548 54654 1584 54660
rect 1548 54651 1554 54654
rect 156 54614 162 54617
rect 126 54608 162 54614
rect 810 54614 816 54617
rect 810 54608 1584 54614
rect 126 54574 138 54608
rect 1572 54574 1584 54608
rect 126 54568 162 54574
rect 156 54565 162 54568
rect 810 54568 1584 54574
rect 810 54565 816 54568
rect 894 54528 900 54531
rect 126 54522 900 54528
rect 1548 54528 1554 54531
rect 1548 54522 1584 54528
rect 126 54488 138 54522
rect 1572 54488 1584 54522
rect 126 54482 900 54488
rect 894 54479 900 54482
rect 1548 54482 1584 54488
rect 1548 54479 1554 54482
rect 156 54442 162 54445
rect 126 54436 162 54442
rect 810 54442 816 54445
rect 810 54436 1584 54442
rect 126 54402 138 54436
rect 1572 54402 1584 54436
rect 126 54396 162 54402
rect 156 54393 162 54396
rect 810 54396 1584 54402
rect 810 54393 816 54396
rect 894 54356 900 54359
rect 126 54350 900 54356
rect 1548 54356 1554 54359
rect 1548 54350 1584 54356
rect 126 54316 138 54350
rect 1572 54316 1584 54350
rect 126 54310 900 54316
rect 894 54307 900 54310
rect 1548 54310 1584 54316
rect 1548 54307 1554 54310
rect 156 54270 162 54273
rect 126 54264 162 54270
rect 810 54270 816 54273
rect 810 54264 1584 54270
rect 126 54230 138 54264
rect 1572 54230 1584 54264
rect 126 54224 162 54230
rect 156 54221 162 54224
rect 810 54224 1584 54230
rect 810 54221 816 54224
rect 894 54184 900 54187
rect 126 54178 900 54184
rect 1548 54184 1554 54187
rect 1548 54178 1584 54184
rect 126 54144 138 54178
rect 1572 54144 1584 54178
rect 126 54138 900 54144
rect 894 54135 900 54138
rect 1548 54138 1584 54144
rect 1548 54135 1554 54138
rect 156 54098 162 54101
rect 126 54092 162 54098
rect 810 54098 816 54101
rect 810 54092 1584 54098
rect 126 54058 138 54092
rect 1572 54058 1584 54092
rect 126 54052 162 54058
rect 156 54049 162 54052
rect 810 54052 1584 54058
rect 810 54049 816 54052
rect 894 54012 900 54015
rect 126 54006 900 54012
rect 1548 54012 1554 54015
rect 1548 54006 1584 54012
rect 126 53972 138 54006
rect 1572 53972 1584 54006
rect 126 53966 900 53972
rect 894 53963 900 53966
rect 1548 53966 1584 53972
rect 1548 53963 1554 53966
rect 156 53926 162 53929
rect 126 53920 162 53926
rect 810 53926 816 53929
rect 810 53920 1584 53926
rect 126 53886 138 53920
rect 1572 53886 1584 53920
rect 126 53880 162 53886
rect 156 53877 162 53880
rect 810 53880 1584 53886
rect 810 53877 816 53880
rect 894 53840 900 53843
rect 126 53834 900 53840
rect 1548 53840 1554 53843
rect 1548 53834 1584 53840
rect 126 53800 138 53834
rect 1572 53800 1584 53834
rect 126 53794 900 53800
rect 894 53791 900 53794
rect 1548 53794 1584 53800
rect 1548 53791 1554 53794
rect 156 53754 162 53757
rect 126 53748 162 53754
rect 810 53754 816 53757
rect 810 53748 1584 53754
rect 126 53714 138 53748
rect 1572 53714 1584 53748
rect 126 53708 162 53714
rect 156 53705 162 53708
rect 810 53708 1584 53714
rect 810 53705 816 53708
rect 894 53668 900 53671
rect 126 53662 900 53668
rect 1548 53668 1554 53671
rect 1548 53662 1584 53668
rect 126 53628 138 53662
rect 1572 53628 1584 53662
rect 126 53622 900 53628
rect 894 53619 900 53622
rect 1548 53622 1584 53628
rect 1548 53619 1554 53622
rect 156 53582 162 53585
rect 126 53576 162 53582
rect 810 53582 816 53585
rect 810 53576 1584 53582
rect 126 53542 138 53576
rect 1572 53542 1584 53576
rect 126 53536 162 53542
rect 156 53533 162 53536
rect 810 53536 1584 53542
rect 810 53533 816 53536
rect 894 53496 900 53499
rect 126 53490 900 53496
rect 1548 53496 1554 53499
rect 1548 53490 1584 53496
rect 126 53456 138 53490
rect 1572 53456 1584 53490
rect 126 53450 900 53456
rect 894 53447 900 53450
rect 1548 53450 1584 53456
rect 1548 53447 1554 53450
rect 156 53410 162 53413
rect 126 53404 162 53410
rect 810 53410 816 53413
rect 810 53404 1584 53410
rect 126 53370 138 53404
rect 1572 53370 1584 53404
rect 126 53364 162 53370
rect 156 53361 162 53364
rect 810 53364 1584 53370
rect 810 53361 816 53364
rect 894 53324 900 53327
rect 126 53318 900 53324
rect 1548 53324 1554 53327
rect 1548 53318 1584 53324
rect 126 53284 138 53318
rect 1572 53284 1584 53318
rect 126 53278 900 53284
rect 894 53275 900 53278
rect 1548 53278 1584 53284
rect 1548 53275 1554 53278
rect 156 53238 162 53241
rect 126 53232 162 53238
rect 810 53238 816 53241
rect 810 53232 1584 53238
rect 126 53198 138 53232
rect 1572 53198 1584 53232
rect 126 53192 162 53198
rect 156 53189 162 53192
rect 810 53192 1584 53198
rect 810 53189 816 53192
rect 894 53152 900 53155
rect 126 53146 900 53152
rect 1548 53152 1554 53155
rect 1548 53146 1584 53152
rect 126 53112 138 53146
rect 1572 53112 1584 53146
rect 126 53106 900 53112
rect 894 53103 900 53106
rect 1548 53106 1584 53112
rect 1548 53103 1554 53106
rect 156 53066 162 53069
rect 126 53060 162 53066
rect 810 53066 816 53069
rect 810 53060 1584 53066
rect 126 53026 138 53060
rect 1572 53026 1584 53060
rect 126 53020 162 53026
rect 156 53017 162 53020
rect 810 53020 1584 53026
rect 810 53017 816 53020
rect 894 52980 900 52983
rect 126 52974 900 52980
rect 1548 52980 1554 52983
rect 1548 52974 1584 52980
rect 126 52940 138 52974
rect 1572 52940 1584 52974
rect 126 52934 900 52940
rect 894 52931 900 52934
rect 1548 52934 1584 52940
rect 1548 52931 1554 52934
rect 156 52894 162 52897
rect 126 52888 162 52894
rect 810 52894 816 52897
rect 810 52888 1584 52894
rect 126 52854 138 52888
rect 1572 52854 1584 52888
rect 126 52848 162 52854
rect 156 52845 162 52848
rect 810 52848 1584 52854
rect 810 52845 816 52848
rect 894 52808 900 52811
rect 126 52802 900 52808
rect 1548 52808 1554 52811
rect 1548 52802 1584 52808
rect 126 52768 138 52802
rect 1572 52768 1584 52802
rect 126 52762 900 52768
rect 894 52759 900 52762
rect 1548 52762 1584 52768
rect 1548 52759 1554 52762
rect 156 52722 162 52725
rect 126 52716 162 52722
rect 810 52722 816 52725
rect 810 52716 1584 52722
rect 126 52682 138 52716
rect 1572 52682 1584 52716
rect 126 52676 162 52682
rect 156 52673 162 52676
rect 810 52676 1584 52682
rect 810 52673 816 52676
rect 894 52636 900 52639
rect 126 52630 900 52636
rect 1548 52636 1554 52639
rect 1548 52630 1584 52636
rect 126 52596 138 52630
rect 1572 52596 1584 52630
rect 126 52590 900 52596
rect 894 52587 900 52590
rect 1548 52590 1584 52596
rect 1548 52587 1554 52590
rect 156 52550 162 52553
rect 126 52544 162 52550
rect 810 52550 816 52553
rect 810 52544 1584 52550
rect 126 52510 138 52544
rect 1572 52510 1584 52544
rect 126 52504 162 52510
rect 156 52501 162 52504
rect 810 52504 1584 52510
rect 810 52501 816 52504
rect 894 52464 900 52467
rect 126 52458 900 52464
rect 1548 52464 1554 52467
rect 1548 52458 1584 52464
rect 126 52424 138 52458
rect 1572 52424 1584 52458
rect 126 52418 900 52424
rect 894 52415 900 52418
rect 1548 52418 1584 52424
rect 1548 52415 1554 52418
rect 156 52378 162 52381
rect 126 52372 162 52378
rect 810 52378 816 52381
rect 810 52372 1584 52378
rect 126 52338 138 52372
rect 1572 52338 1584 52372
rect 126 52332 162 52338
rect 156 52329 162 52332
rect 810 52332 1584 52338
rect 810 52329 816 52332
rect 894 52292 900 52295
rect 126 52286 900 52292
rect 1548 52292 1554 52295
rect 1548 52286 1584 52292
rect 126 52252 138 52286
rect 1572 52252 1584 52286
rect 126 52246 900 52252
rect 894 52243 900 52246
rect 1548 52246 1584 52252
rect 1548 52243 1554 52246
rect 156 52206 162 52209
rect 126 52200 162 52206
rect 810 52206 816 52209
rect 810 52200 1584 52206
rect 126 52166 138 52200
rect 1572 52166 1584 52200
rect 126 52160 162 52166
rect 156 52157 162 52160
rect 810 52160 1584 52166
rect 810 52157 816 52160
rect 894 52120 900 52123
rect 126 52114 900 52120
rect 1548 52120 1554 52123
rect 1548 52114 1584 52120
rect 126 52080 138 52114
rect 1572 52080 1584 52114
rect 126 52074 900 52080
rect 894 52071 900 52074
rect 1548 52074 1584 52080
rect 1548 52071 1554 52074
rect 156 52034 162 52037
rect 126 52028 162 52034
rect 810 52034 816 52037
rect 810 52028 1584 52034
rect 126 51994 138 52028
rect 1572 51994 1584 52028
rect 126 51988 162 51994
rect 156 51985 162 51988
rect 810 51988 1584 51994
rect 810 51985 816 51988
rect 894 51948 900 51951
rect 126 51942 900 51948
rect 1548 51948 1554 51951
rect 1548 51942 1584 51948
rect 126 51908 138 51942
rect 1572 51908 1584 51942
rect 126 51902 900 51908
rect 894 51899 900 51902
rect 1548 51902 1584 51908
rect 1548 51899 1554 51902
rect 156 51862 162 51865
rect 126 51856 162 51862
rect 810 51862 816 51865
rect 810 51856 1584 51862
rect 126 51822 138 51856
rect 1572 51822 1584 51856
rect 126 51816 162 51822
rect 156 51813 162 51816
rect 810 51816 1584 51822
rect 810 51813 816 51816
rect 894 51776 900 51779
rect 126 51770 900 51776
rect 1548 51776 1554 51779
rect 1548 51770 1584 51776
rect 126 51736 138 51770
rect 1572 51736 1584 51770
rect 126 51730 900 51736
rect 894 51727 900 51730
rect 1548 51730 1584 51736
rect 1548 51727 1554 51730
rect 156 51690 162 51693
rect 126 51684 162 51690
rect 810 51690 816 51693
rect 810 51684 1584 51690
rect 126 51650 138 51684
rect 1572 51650 1584 51684
rect 126 51644 162 51650
rect 156 51641 162 51644
rect 810 51644 1584 51650
rect 810 51641 816 51644
rect 894 51604 900 51607
rect 126 51598 900 51604
rect 1548 51604 1554 51607
rect 1548 51598 1584 51604
rect 126 51564 138 51598
rect 1572 51564 1584 51598
rect 126 51558 900 51564
rect 894 51555 900 51558
rect 1548 51558 1584 51564
rect 1548 51555 1554 51558
rect 156 51518 162 51521
rect 126 51512 162 51518
rect 810 51518 816 51521
rect 810 51512 1584 51518
rect 126 51478 138 51512
rect 1572 51478 1584 51512
rect 126 51472 162 51478
rect 156 51469 162 51472
rect 810 51472 1584 51478
rect 810 51469 816 51472
rect 894 51432 900 51435
rect 126 51426 900 51432
rect 1548 51432 1554 51435
rect 1548 51426 1584 51432
rect 126 51392 138 51426
rect 1572 51392 1584 51426
rect 126 51386 900 51392
rect 894 51383 900 51386
rect 1548 51386 1584 51392
rect 1548 51383 1554 51386
rect 156 51346 162 51349
rect 126 51340 162 51346
rect 810 51346 816 51349
rect 810 51340 1584 51346
rect 126 51306 138 51340
rect 1572 51306 1584 51340
rect 126 51300 162 51306
rect 156 51297 162 51300
rect 810 51300 1584 51306
rect 810 51297 816 51300
rect 894 51260 900 51263
rect 126 51254 900 51260
rect 1548 51260 1554 51263
rect 1548 51254 1584 51260
rect 126 51220 138 51254
rect 1572 51220 1584 51254
rect 126 51214 900 51220
rect 894 51211 900 51214
rect 1548 51214 1584 51220
rect 1548 51211 1554 51214
rect 156 51174 162 51177
rect 126 51168 162 51174
rect 810 51174 816 51177
rect 810 51168 1584 51174
rect 126 51134 138 51168
rect 1572 51134 1584 51168
rect 126 51128 162 51134
rect 156 51125 162 51128
rect 810 51128 1584 51134
rect 810 51125 816 51128
rect 894 51088 900 51091
rect 126 51082 900 51088
rect 1548 51088 1554 51091
rect 1548 51082 1584 51088
rect 126 51048 138 51082
rect 1572 51048 1584 51082
rect 126 51042 900 51048
rect 894 51039 900 51042
rect 1548 51042 1584 51048
rect 1548 51039 1554 51042
rect 156 51002 162 51005
rect 126 50996 162 51002
rect 810 51002 816 51005
rect 810 50996 1584 51002
rect 126 50962 138 50996
rect 1572 50962 1584 50996
rect 126 50956 162 50962
rect 156 50953 162 50956
rect 810 50956 1584 50962
rect 810 50953 816 50956
rect 894 50916 900 50919
rect 126 50910 900 50916
rect 1548 50916 1554 50919
rect 1548 50910 1584 50916
rect 126 50876 138 50910
rect 1572 50876 1584 50910
rect 126 50870 900 50876
rect 894 50867 900 50870
rect 1548 50870 1584 50876
rect 1548 50867 1554 50870
rect 156 50830 162 50833
rect 126 50824 162 50830
rect 810 50830 816 50833
rect 810 50824 1584 50830
rect 126 50790 138 50824
rect 1572 50790 1584 50824
rect 126 50784 162 50790
rect 156 50781 162 50784
rect 810 50784 1584 50790
rect 810 50781 816 50784
rect 894 50744 900 50747
rect 126 50738 900 50744
rect 1548 50744 1554 50747
rect 1548 50738 1584 50744
rect 126 50704 138 50738
rect 1572 50704 1584 50738
rect 126 50698 900 50704
rect 894 50695 900 50698
rect 1548 50698 1584 50704
rect 1548 50695 1554 50698
rect 156 50658 162 50661
rect 126 50652 162 50658
rect 810 50658 816 50661
rect 810 50652 1584 50658
rect 126 50618 138 50652
rect 1572 50618 1584 50652
rect 126 50612 162 50618
rect 156 50609 162 50612
rect 810 50612 1584 50618
rect 810 50609 816 50612
rect 894 50572 900 50575
rect 126 50566 900 50572
rect 1548 50572 1554 50575
rect 1548 50566 1584 50572
rect 126 50532 138 50566
rect 1572 50532 1584 50566
rect 126 50526 900 50532
rect 894 50523 900 50526
rect 1548 50526 1584 50532
rect 1548 50523 1554 50526
rect 156 50486 162 50489
rect 126 50480 162 50486
rect 810 50486 816 50489
rect 810 50480 1584 50486
rect 126 50446 138 50480
rect 1572 50446 1584 50480
rect 126 50440 162 50446
rect 156 50437 162 50440
rect 810 50440 1584 50446
rect 810 50437 816 50440
rect 894 50400 900 50403
rect 126 50394 900 50400
rect 1548 50400 1554 50403
rect 1548 50394 1584 50400
rect 126 50360 138 50394
rect 1572 50360 1584 50394
rect 126 50354 900 50360
rect 894 50351 900 50354
rect 1548 50354 1584 50360
rect 1548 50351 1554 50354
rect 156 50314 162 50317
rect 126 50308 162 50314
rect 810 50314 816 50317
rect 810 50308 1584 50314
rect 126 50274 138 50308
rect 1572 50274 1584 50308
rect 126 50268 162 50274
rect 156 50265 162 50268
rect 810 50268 1584 50274
rect 810 50265 816 50268
rect 894 50228 900 50231
rect 126 50222 900 50228
rect 1548 50228 1554 50231
rect 1548 50222 1584 50228
rect 126 50188 138 50222
rect 1572 50188 1584 50222
rect 126 50182 900 50188
rect 894 50179 900 50182
rect 1548 50182 1584 50188
rect 1548 50179 1554 50182
rect 156 50142 162 50145
rect 126 50136 162 50142
rect 810 50142 816 50145
rect 810 50136 1584 50142
rect 126 50102 138 50136
rect 1572 50102 1584 50136
rect 126 50096 162 50102
rect 156 50093 162 50096
rect 810 50096 1584 50102
rect 810 50093 816 50096
rect 894 50056 900 50059
rect 126 50050 900 50056
rect 1548 50056 1554 50059
rect 1548 50050 1584 50056
rect 126 50016 138 50050
rect 1572 50016 1584 50050
rect 126 50010 900 50016
rect 894 50007 900 50010
rect 1548 50010 1584 50016
rect 1548 50007 1554 50010
rect 156 49970 162 49973
rect 126 49964 162 49970
rect 810 49970 816 49973
rect 810 49964 1584 49970
rect 126 49930 138 49964
rect 1572 49930 1584 49964
rect 126 49924 162 49930
rect 156 49921 162 49924
rect 810 49924 1584 49930
rect 810 49921 816 49924
rect 894 49884 900 49887
rect 126 49878 900 49884
rect 1548 49884 1554 49887
rect 1548 49878 1584 49884
rect 126 49844 138 49878
rect 1572 49844 1584 49878
rect 126 49838 900 49844
rect 894 49835 900 49838
rect 1548 49838 1584 49844
rect 1548 49835 1554 49838
rect 156 49798 162 49801
rect 126 49792 162 49798
rect 810 49798 816 49801
rect 810 49792 1584 49798
rect 126 49758 138 49792
rect 1572 49758 1584 49792
rect 126 49752 162 49758
rect 156 49749 162 49752
rect 810 49752 1584 49758
rect 810 49749 816 49752
rect 894 49712 900 49715
rect 126 49706 900 49712
rect 1548 49712 1554 49715
rect 1548 49706 1584 49712
rect 126 49672 138 49706
rect 1572 49672 1584 49706
rect 126 49666 900 49672
rect 894 49663 900 49666
rect 1548 49666 1584 49672
rect 1548 49663 1554 49666
rect 156 49626 162 49629
rect 126 49620 162 49626
rect 810 49626 816 49629
rect 810 49620 1584 49626
rect 126 49586 138 49620
rect 1572 49586 1584 49620
rect 126 49580 162 49586
rect 156 49577 162 49580
rect 810 49580 1584 49586
rect 810 49577 816 49580
rect 894 49540 900 49543
rect 126 49534 900 49540
rect 1548 49540 1554 49543
rect 1548 49534 1584 49540
rect 126 49500 138 49534
rect 1572 49500 1584 49534
rect 126 49494 900 49500
rect 894 49491 900 49494
rect 1548 49494 1584 49500
rect 1548 49491 1554 49494
rect 156 49454 162 49457
rect 126 49448 162 49454
rect 810 49454 816 49457
rect 810 49448 1584 49454
rect 126 49414 138 49448
rect 1572 49414 1584 49448
rect 126 49408 162 49414
rect 156 49405 162 49408
rect 810 49408 1584 49414
rect 810 49405 816 49408
rect 894 49368 900 49371
rect 126 49362 900 49368
rect 1548 49368 1554 49371
rect 1548 49362 1584 49368
rect 126 49328 138 49362
rect 1572 49328 1584 49362
rect 126 49322 900 49328
rect 894 49319 900 49322
rect 1548 49322 1584 49328
rect 1548 49319 1554 49322
rect 156 49282 162 49285
rect 126 49276 162 49282
rect 810 49282 816 49285
rect 810 49276 1584 49282
rect 126 49242 138 49276
rect 1572 49242 1584 49276
rect 126 49236 162 49242
rect 156 49233 162 49236
rect 810 49236 1584 49242
rect 810 49233 816 49236
rect 894 49196 900 49199
rect 126 49190 900 49196
rect 1548 49196 1554 49199
rect 1548 49190 1584 49196
rect 126 49156 138 49190
rect 1572 49156 1584 49190
rect 126 49150 900 49156
rect 894 49147 900 49150
rect 1548 49150 1584 49156
rect 1548 49147 1554 49150
rect 156 49110 162 49113
rect 126 49104 162 49110
rect 810 49110 816 49113
rect 810 49104 1584 49110
rect 126 49070 138 49104
rect 1572 49070 1584 49104
rect 126 49064 162 49070
rect 156 49061 162 49064
rect 810 49064 1584 49070
rect 810 49061 816 49064
rect 894 49024 900 49027
rect 126 49018 900 49024
rect 1548 49024 1554 49027
rect 1548 49018 1584 49024
rect 126 48984 138 49018
rect 1572 48984 1584 49018
rect 126 48978 900 48984
rect 894 48975 900 48978
rect 1548 48978 1584 48984
rect 1548 48975 1554 48978
rect 156 48938 162 48941
rect 126 48932 162 48938
rect 810 48938 816 48941
rect 810 48932 1584 48938
rect 126 48898 138 48932
rect 1572 48898 1584 48932
rect 126 48892 162 48898
rect 156 48889 162 48892
rect 810 48892 1584 48898
rect 810 48889 816 48892
rect 894 48852 900 48855
rect 126 48846 900 48852
rect 1548 48852 1554 48855
rect 1548 48846 1584 48852
rect 126 48812 138 48846
rect 1572 48812 1584 48846
rect 126 48806 900 48812
rect 894 48803 900 48806
rect 1548 48806 1584 48812
rect 1548 48803 1554 48806
rect 156 48766 162 48769
rect 126 48760 162 48766
rect 810 48766 816 48769
rect 810 48760 1584 48766
rect 126 48726 138 48760
rect 1572 48726 1584 48760
rect 126 48720 162 48726
rect 156 48717 162 48720
rect 810 48720 1584 48726
rect 810 48717 816 48720
rect 894 48680 900 48683
rect 126 48674 900 48680
rect 1548 48680 1554 48683
rect 1548 48674 1584 48680
rect 126 48640 138 48674
rect 1572 48640 1584 48674
rect 126 48634 900 48640
rect 894 48631 900 48634
rect 1548 48634 1584 48640
rect 1548 48631 1554 48634
rect 156 48594 162 48597
rect 126 48588 162 48594
rect 810 48594 816 48597
rect 810 48588 1584 48594
rect 126 48554 138 48588
rect 1572 48554 1584 48588
rect 126 48548 162 48554
rect 156 48545 162 48548
rect 810 48548 1584 48554
rect 810 48545 816 48548
rect 894 48508 900 48511
rect 126 48502 900 48508
rect 1548 48508 1554 48511
rect 1548 48502 1584 48508
rect 126 48468 138 48502
rect 1572 48468 1584 48502
rect 126 48462 900 48468
rect 894 48459 900 48462
rect 1548 48462 1584 48468
rect 1548 48459 1554 48462
rect 156 48422 162 48425
rect 126 48416 162 48422
rect 810 48422 816 48425
rect 810 48416 1584 48422
rect 126 48382 138 48416
rect 1572 48382 1584 48416
rect 126 48376 162 48382
rect 156 48373 162 48376
rect 810 48376 1584 48382
rect 810 48373 816 48376
rect 894 48336 900 48339
rect 126 48330 900 48336
rect 1548 48336 1554 48339
rect 1548 48330 1584 48336
rect 126 48296 138 48330
rect 1572 48296 1584 48330
rect 126 48290 900 48296
rect 894 48287 900 48290
rect 1548 48290 1584 48296
rect 1548 48287 1554 48290
rect 156 48250 162 48253
rect 126 48244 162 48250
rect 810 48250 816 48253
rect 810 48244 1584 48250
rect 126 48210 138 48244
rect 1572 48210 1584 48244
rect 126 48204 162 48210
rect 156 48201 162 48204
rect 810 48204 1584 48210
rect 810 48201 816 48204
rect 894 48164 900 48167
rect 126 48158 900 48164
rect 1548 48164 1554 48167
rect 1548 48158 1584 48164
rect 126 48124 138 48158
rect 1572 48124 1584 48158
rect 126 48118 900 48124
rect 894 48115 900 48118
rect 1548 48118 1584 48124
rect 1548 48115 1554 48118
rect 156 48078 162 48081
rect 126 48072 162 48078
rect 810 48078 816 48081
rect 810 48072 1584 48078
rect 126 48038 138 48072
rect 1572 48038 1584 48072
rect 126 48032 162 48038
rect 156 48029 162 48032
rect 810 48032 1584 48038
rect 810 48029 816 48032
rect 894 47992 900 47995
rect 126 47986 900 47992
rect 1548 47992 1554 47995
rect 1548 47986 1584 47992
rect 126 47952 138 47986
rect 1572 47952 1584 47986
rect 126 47946 900 47952
rect 894 47943 900 47946
rect 1548 47946 1584 47952
rect 1548 47943 1554 47946
rect 156 47906 162 47909
rect 126 47900 162 47906
rect 810 47906 816 47909
rect 810 47900 1584 47906
rect 126 47866 138 47900
rect 1572 47866 1584 47900
rect 126 47860 162 47866
rect 156 47857 162 47860
rect 810 47860 1584 47866
rect 810 47857 816 47860
rect 894 47820 900 47823
rect 126 47814 900 47820
rect 1548 47820 1554 47823
rect 1548 47814 1584 47820
rect 126 47780 138 47814
rect 1572 47780 1584 47814
rect 126 47774 900 47780
rect 894 47771 900 47774
rect 1548 47774 1584 47780
rect 1548 47771 1554 47774
rect 156 47734 162 47737
rect 126 47728 162 47734
rect 810 47734 816 47737
rect 810 47728 1584 47734
rect 126 47694 138 47728
rect 1572 47694 1584 47728
rect 126 47688 162 47694
rect 156 47685 162 47688
rect 810 47688 1584 47694
rect 810 47685 816 47688
rect 894 47648 900 47651
rect 126 47642 900 47648
rect 1548 47648 1554 47651
rect 1548 47642 1584 47648
rect 126 47608 138 47642
rect 1572 47608 1584 47642
rect 126 47602 900 47608
rect 894 47599 900 47602
rect 1548 47602 1584 47608
rect 1548 47599 1554 47602
rect 156 47562 162 47565
rect 126 47556 162 47562
rect 810 47562 816 47565
rect 810 47556 1584 47562
rect 126 47522 138 47556
rect 1572 47522 1584 47556
rect 126 47516 162 47522
rect 156 47513 162 47516
rect 810 47516 1584 47522
rect 810 47513 816 47516
rect 894 47476 900 47479
rect 126 47470 900 47476
rect 1548 47476 1554 47479
rect 1548 47470 1584 47476
rect 126 47436 138 47470
rect 1572 47436 1584 47470
rect 126 47430 900 47436
rect 894 47427 900 47430
rect 1548 47430 1584 47436
rect 1548 47427 1554 47430
rect 156 47390 162 47393
rect 126 47384 162 47390
rect 810 47390 816 47393
rect 810 47384 1584 47390
rect 126 47350 138 47384
rect 1572 47350 1584 47384
rect 126 47344 162 47350
rect 156 47341 162 47344
rect 810 47344 1584 47350
rect 810 47341 816 47344
rect 894 47304 900 47307
rect 126 47298 900 47304
rect 1548 47304 1554 47307
rect 1548 47298 1584 47304
rect 126 47264 138 47298
rect 1572 47264 1584 47298
rect 126 47258 900 47264
rect 894 47255 900 47258
rect 1548 47258 1584 47264
rect 1548 47255 1554 47258
rect 156 47218 162 47221
rect 126 47212 162 47218
rect 810 47218 816 47221
rect 810 47212 1584 47218
rect 126 47178 138 47212
rect 1572 47178 1584 47212
rect 126 47172 162 47178
rect 156 47169 162 47172
rect 810 47172 1584 47178
rect 810 47169 816 47172
rect 894 47132 900 47135
rect 126 47126 900 47132
rect 1548 47132 1554 47135
rect 1548 47126 1584 47132
rect 126 47092 138 47126
rect 1572 47092 1584 47126
rect 126 47086 900 47092
rect 894 47083 900 47086
rect 1548 47086 1584 47092
rect 1548 47083 1554 47086
rect 156 47046 162 47049
rect 126 47040 162 47046
rect 810 47046 816 47049
rect 810 47040 1584 47046
rect 126 47006 138 47040
rect 1572 47006 1584 47040
rect 126 47000 162 47006
rect 156 46997 162 47000
rect 810 47000 1584 47006
rect 810 46997 816 47000
rect 894 46960 900 46963
rect 126 46954 900 46960
rect 1548 46960 1554 46963
rect 1548 46954 1584 46960
rect 126 46920 138 46954
rect 1572 46920 1584 46954
rect 126 46914 900 46920
rect 894 46911 900 46914
rect 1548 46914 1584 46920
rect 1548 46911 1554 46914
rect 156 46874 162 46877
rect 126 46868 162 46874
rect 810 46874 816 46877
rect 810 46868 1584 46874
rect 126 46834 138 46868
rect 1572 46834 1584 46868
rect 126 46828 162 46834
rect 156 46825 162 46828
rect 810 46828 1584 46834
rect 810 46825 816 46828
rect 894 46788 900 46791
rect 126 46782 900 46788
rect 1548 46788 1554 46791
rect 1548 46782 1584 46788
rect 126 46748 138 46782
rect 1572 46748 1584 46782
rect 126 46742 900 46748
rect 894 46739 900 46742
rect 1548 46742 1584 46748
rect 1548 46739 1554 46742
rect 156 46702 162 46705
rect 126 46696 162 46702
rect 810 46702 816 46705
rect 810 46696 1584 46702
rect 126 46662 138 46696
rect 1572 46662 1584 46696
rect 126 46656 162 46662
rect 156 46653 162 46656
rect 810 46656 1584 46662
rect 810 46653 816 46656
rect 894 46616 900 46619
rect 126 46610 900 46616
rect 1548 46616 1554 46619
rect 1548 46610 1584 46616
rect 126 46576 138 46610
rect 1572 46576 1584 46610
rect 126 46570 900 46576
rect 894 46567 900 46570
rect 1548 46570 1584 46576
rect 1548 46567 1554 46570
rect 156 46530 162 46533
rect 126 46524 162 46530
rect 810 46530 816 46533
rect 810 46524 1584 46530
rect 126 46490 138 46524
rect 1572 46490 1584 46524
rect 126 46484 162 46490
rect 156 46481 162 46484
rect 810 46484 1584 46490
rect 810 46481 816 46484
rect 894 46444 900 46447
rect 126 46438 900 46444
rect 1548 46444 1554 46447
rect 1548 46438 1584 46444
rect 126 46404 138 46438
rect 1572 46404 1584 46438
rect 126 46398 900 46404
rect 894 46395 900 46398
rect 1548 46398 1584 46404
rect 1548 46395 1554 46398
rect 156 46358 162 46361
rect 126 46352 162 46358
rect 810 46358 816 46361
rect 810 46352 1584 46358
rect 126 46318 138 46352
rect 1572 46318 1584 46352
rect 126 46312 162 46318
rect 156 46309 162 46312
rect 810 46312 1584 46318
rect 810 46309 816 46312
rect 894 46272 900 46275
rect 126 46266 900 46272
rect 1548 46272 1554 46275
rect 1548 46266 1584 46272
rect 126 46232 138 46266
rect 1572 46232 1584 46266
rect 126 46226 900 46232
rect 894 46223 900 46226
rect 1548 46226 1584 46232
rect 1548 46223 1554 46226
rect 156 46186 162 46189
rect 126 46180 162 46186
rect 810 46186 816 46189
rect 810 46180 1584 46186
rect 126 46146 138 46180
rect 1572 46146 1584 46180
rect 126 46140 162 46146
rect 156 46137 162 46140
rect 810 46140 1584 46146
rect 810 46137 816 46140
rect 894 46100 900 46103
rect 126 46094 900 46100
rect 1548 46100 1554 46103
rect 1548 46094 1584 46100
rect 126 46060 138 46094
rect 1572 46060 1584 46094
rect 126 46054 900 46060
rect 894 46051 900 46054
rect 1548 46054 1584 46060
rect 1548 46051 1554 46054
rect 156 46014 162 46017
rect 126 46008 162 46014
rect 810 46014 816 46017
rect 810 46008 1584 46014
rect 126 45974 138 46008
rect 1572 45974 1584 46008
rect 126 45968 162 45974
rect 156 45965 162 45968
rect 810 45968 1584 45974
rect 810 45965 816 45968
rect 894 45928 900 45931
rect 126 45922 900 45928
rect 1548 45928 1554 45931
rect 1548 45922 1584 45928
rect 126 45888 138 45922
rect 1572 45888 1584 45922
rect 126 45882 900 45888
rect 894 45879 900 45882
rect 1548 45882 1584 45888
rect 1548 45879 1554 45882
rect 156 45842 162 45845
rect 126 45836 162 45842
rect 810 45842 816 45845
rect 810 45836 1584 45842
rect 126 45802 138 45836
rect 1572 45802 1584 45836
rect 126 45796 162 45802
rect 156 45793 162 45796
rect 810 45796 1584 45802
rect 810 45793 816 45796
rect 894 45756 900 45759
rect 126 45750 900 45756
rect 1548 45756 1554 45759
rect 1548 45750 1584 45756
rect 126 45716 138 45750
rect 1572 45716 1584 45750
rect 126 45710 900 45716
rect 894 45707 900 45710
rect 1548 45710 1584 45716
rect 1548 45707 1554 45710
rect 156 45670 162 45673
rect 126 45664 162 45670
rect 810 45670 816 45673
rect 810 45664 1584 45670
rect 126 45630 138 45664
rect 1572 45630 1584 45664
rect 126 45624 162 45630
rect 156 45621 162 45624
rect 810 45624 1584 45630
rect 810 45621 816 45624
rect 894 45584 900 45587
rect 126 45578 900 45584
rect 1548 45584 1554 45587
rect 1548 45578 1584 45584
rect 126 45544 138 45578
rect 1572 45544 1584 45578
rect 126 45538 900 45544
rect 894 45535 900 45538
rect 1548 45538 1584 45544
rect 1548 45535 1554 45538
rect 156 45498 162 45501
rect 126 45492 162 45498
rect 810 45498 816 45501
rect 810 45492 1584 45498
rect 126 45458 138 45492
rect 1572 45458 1584 45492
rect 126 45452 162 45458
rect 156 45449 162 45452
rect 810 45452 1584 45458
rect 810 45449 816 45452
rect 894 45412 900 45415
rect 126 45406 900 45412
rect 1548 45412 1554 45415
rect 1548 45406 1584 45412
rect 126 45372 138 45406
rect 1572 45372 1584 45406
rect 126 45366 900 45372
rect 894 45363 900 45366
rect 1548 45366 1584 45372
rect 1548 45363 1554 45366
rect 156 45326 162 45329
rect 126 45320 162 45326
rect 810 45326 816 45329
rect 810 45320 1584 45326
rect 126 45286 138 45320
rect 1572 45286 1584 45320
rect 126 45280 162 45286
rect 156 45277 162 45280
rect 810 45280 1584 45286
rect 810 45277 816 45280
rect 894 45240 900 45243
rect 126 45234 900 45240
rect 1548 45240 1554 45243
rect 1548 45234 1584 45240
rect 126 45200 138 45234
rect 1572 45200 1584 45234
rect 126 45194 900 45200
rect 894 45191 900 45194
rect 1548 45194 1584 45200
rect 1548 45191 1554 45194
rect 156 45154 162 45157
rect 126 45148 162 45154
rect 810 45154 816 45157
rect 810 45148 1584 45154
rect 126 45114 138 45148
rect 1572 45114 1584 45148
rect 126 45108 162 45114
rect 156 45105 162 45108
rect 810 45108 1584 45114
rect 810 45105 816 45108
rect 894 45068 900 45071
rect 126 45062 900 45068
rect 1548 45068 1554 45071
rect 1548 45062 1584 45068
rect 126 45028 138 45062
rect 1572 45028 1584 45062
rect 126 45022 900 45028
rect 894 45019 900 45022
rect 1548 45022 1584 45028
rect 1548 45019 1554 45022
rect 156 44982 162 44985
rect 126 44976 162 44982
rect 810 44982 816 44985
rect 810 44976 1584 44982
rect 126 44942 138 44976
rect 1572 44942 1584 44976
rect 126 44936 162 44942
rect 156 44933 162 44936
rect 810 44936 1584 44942
rect 810 44933 816 44936
rect 894 44896 900 44899
rect 126 44890 900 44896
rect 1548 44896 1554 44899
rect 1548 44890 1584 44896
rect 126 44856 138 44890
rect 1572 44856 1584 44890
rect 126 44850 900 44856
rect 894 44847 900 44850
rect 1548 44850 1584 44856
rect 1548 44847 1554 44850
rect 156 44810 162 44813
rect 126 44804 162 44810
rect 810 44810 816 44813
rect 810 44804 1584 44810
rect 126 44770 138 44804
rect 1572 44770 1584 44804
rect 126 44764 162 44770
rect 156 44761 162 44764
rect 810 44764 1584 44770
rect 810 44761 816 44764
rect 894 44724 900 44727
rect 126 44718 900 44724
rect 1548 44724 1554 44727
rect 1548 44718 1584 44724
rect 126 44684 138 44718
rect 1572 44684 1584 44718
rect 126 44678 900 44684
rect 894 44675 900 44678
rect 1548 44678 1584 44684
rect 1548 44675 1554 44678
rect 156 44638 162 44641
rect 126 44632 162 44638
rect 810 44638 816 44641
rect 810 44632 1584 44638
rect 126 44598 138 44632
rect 1572 44598 1584 44632
rect 126 44592 162 44598
rect 156 44589 162 44592
rect 810 44592 1584 44598
rect 810 44589 816 44592
rect 894 44552 900 44555
rect 126 44546 900 44552
rect 1548 44552 1554 44555
rect 1548 44546 1584 44552
rect 126 44512 138 44546
rect 1572 44512 1584 44546
rect 126 44506 900 44512
rect 894 44503 900 44506
rect 1548 44506 1584 44512
rect 1548 44503 1554 44506
rect 156 44466 162 44469
rect 126 44460 162 44466
rect 810 44466 816 44469
rect 810 44460 1584 44466
rect 126 44426 138 44460
rect 1572 44426 1584 44460
rect 126 44420 162 44426
rect 156 44417 162 44420
rect 810 44420 1584 44426
rect 810 44417 816 44420
rect 894 44380 900 44383
rect 126 44374 900 44380
rect 1548 44380 1554 44383
rect 1548 44374 1584 44380
rect 126 44340 138 44374
rect 1572 44340 1584 44374
rect 126 44334 900 44340
rect 894 44331 900 44334
rect 1548 44334 1584 44340
rect 1548 44331 1554 44334
rect 156 44294 162 44297
rect 126 44288 162 44294
rect 810 44294 816 44297
rect 810 44288 1584 44294
rect 126 44254 138 44288
rect 1572 44254 1584 44288
rect 126 44248 162 44254
rect 156 44245 162 44248
rect 810 44248 1584 44254
rect 810 44245 816 44248
rect 894 44208 900 44211
rect 126 44202 900 44208
rect 1548 44208 1554 44211
rect 1548 44202 1584 44208
rect 126 44168 138 44202
rect 1572 44168 1584 44202
rect 126 44162 900 44168
rect 894 44159 900 44162
rect 1548 44162 1584 44168
rect 1548 44159 1554 44162
rect 156 44122 162 44125
rect 126 44116 162 44122
rect 810 44122 816 44125
rect 810 44116 1584 44122
rect 126 44082 138 44116
rect 1572 44082 1584 44116
rect 126 44076 162 44082
rect 156 44073 162 44076
rect 810 44076 1584 44082
rect 810 44073 816 44076
rect 894 44036 900 44039
rect 126 44030 900 44036
rect 1548 44036 1554 44039
rect 1548 44030 1584 44036
rect 126 43996 138 44030
rect 1572 43996 1584 44030
rect 126 43990 900 43996
rect 894 43987 900 43990
rect 1548 43990 1584 43996
rect 1548 43987 1554 43990
rect 156 43950 162 43953
rect 126 43944 162 43950
rect 810 43950 816 43953
rect 810 43944 1584 43950
rect 126 43910 138 43944
rect 1572 43910 1584 43944
rect 126 43904 162 43910
rect 156 43901 162 43904
rect 810 43904 1584 43910
rect 810 43901 816 43904
rect 894 43864 900 43867
rect 126 43858 900 43864
rect 1548 43864 1554 43867
rect 1548 43858 1584 43864
rect 126 43824 138 43858
rect 1572 43824 1584 43858
rect 126 43818 900 43824
rect 894 43815 900 43818
rect 1548 43818 1584 43824
rect 1548 43815 1554 43818
rect 156 43778 162 43781
rect 126 43772 162 43778
rect 810 43778 816 43781
rect 810 43772 1584 43778
rect 126 43738 138 43772
rect 1572 43738 1584 43772
rect 126 43732 162 43738
rect 156 43729 162 43732
rect 810 43732 1584 43738
rect 810 43729 816 43732
rect 894 43692 900 43695
rect 126 43686 900 43692
rect 1548 43692 1554 43695
rect 1548 43686 1584 43692
rect 126 43652 138 43686
rect 1572 43652 1584 43686
rect 126 43646 900 43652
rect 894 43643 900 43646
rect 1548 43646 1584 43652
rect 1548 43643 1554 43646
rect 156 43606 162 43609
rect 126 43600 162 43606
rect 810 43606 816 43609
rect 810 43600 1584 43606
rect 126 43566 138 43600
rect 1572 43566 1584 43600
rect 126 43560 162 43566
rect 156 43557 162 43560
rect 810 43560 1584 43566
rect 810 43557 816 43560
rect 894 43520 900 43523
rect 126 43514 900 43520
rect 1548 43520 1554 43523
rect 1548 43514 1584 43520
rect 126 43480 138 43514
rect 1572 43480 1584 43514
rect 126 43474 900 43480
rect 894 43471 900 43474
rect 1548 43474 1584 43480
rect 1548 43471 1554 43474
rect 156 43434 162 43437
rect 126 43428 162 43434
rect 810 43434 816 43437
rect 810 43428 1584 43434
rect 126 43394 138 43428
rect 1572 43394 1584 43428
rect 126 43388 162 43394
rect 156 43385 162 43388
rect 810 43388 1584 43394
rect 810 43385 816 43388
rect 894 43348 900 43351
rect 126 43342 900 43348
rect 1548 43348 1554 43351
rect 1548 43342 1584 43348
rect 126 43308 138 43342
rect 1572 43308 1584 43342
rect 126 43302 900 43308
rect 894 43299 900 43302
rect 1548 43302 1584 43308
rect 1548 43299 1554 43302
rect 156 43262 162 43265
rect 126 43256 162 43262
rect 810 43262 816 43265
rect 810 43256 1584 43262
rect 126 43222 138 43256
rect 1572 43222 1584 43256
rect 126 43216 162 43222
rect 156 43213 162 43216
rect 810 43216 1584 43222
rect 810 43213 816 43216
rect 894 43176 900 43179
rect 126 43170 900 43176
rect 1548 43176 1554 43179
rect 1548 43170 1584 43176
rect 126 43136 138 43170
rect 1572 43136 1584 43170
rect 126 43130 900 43136
rect 894 43127 900 43130
rect 1548 43130 1584 43136
rect 1548 43127 1554 43130
rect 156 43090 162 43093
rect 126 43084 162 43090
rect 810 43090 816 43093
rect 810 43084 1584 43090
rect 126 43050 138 43084
rect 1572 43050 1584 43084
rect 126 43044 162 43050
rect 156 43041 162 43044
rect 810 43044 1584 43050
rect 810 43041 816 43044
rect 894 43004 900 43007
rect 126 42998 900 43004
rect 1548 43004 1554 43007
rect 1548 42998 1584 43004
rect 126 42964 138 42998
rect 1572 42964 1584 42998
rect 126 42958 900 42964
rect 894 42955 900 42958
rect 1548 42958 1584 42964
rect 1548 42955 1554 42958
rect 156 42918 162 42921
rect 126 42912 162 42918
rect 810 42918 816 42921
rect 810 42912 1584 42918
rect 126 42878 138 42912
rect 1572 42878 1584 42912
rect 126 42872 162 42878
rect 156 42869 162 42872
rect 810 42872 1584 42878
rect 810 42869 816 42872
rect 894 42832 900 42835
rect 126 42826 900 42832
rect 1548 42832 1554 42835
rect 1548 42826 1584 42832
rect 126 42792 138 42826
rect 1572 42792 1584 42826
rect 126 42786 900 42792
rect 894 42783 900 42786
rect 1548 42786 1584 42792
rect 1548 42783 1554 42786
rect 156 42746 162 42749
rect 126 42740 162 42746
rect 810 42746 816 42749
rect 810 42740 1584 42746
rect 126 42706 138 42740
rect 1572 42706 1584 42740
rect 126 42700 162 42706
rect 156 42697 162 42700
rect 810 42700 1584 42706
rect 810 42697 816 42700
rect 894 42660 900 42663
rect 126 42654 900 42660
rect 1548 42660 1554 42663
rect 1548 42654 1584 42660
rect 126 42620 138 42654
rect 1572 42620 1584 42654
rect 126 42614 900 42620
rect 894 42611 900 42614
rect 1548 42614 1584 42620
rect 1548 42611 1554 42614
rect 156 42574 162 42577
rect 126 42568 162 42574
rect 810 42574 816 42577
rect 810 42568 1584 42574
rect 126 42534 138 42568
rect 1572 42534 1584 42568
rect 126 42528 162 42534
rect 156 42525 162 42528
rect 810 42528 1584 42534
rect 810 42525 816 42528
rect 894 42488 900 42491
rect 126 42482 900 42488
rect 1548 42488 1554 42491
rect 1548 42482 1584 42488
rect 126 42448 138 42482
rect 1572 42448 1584 42482
rect 126 42442 900 42448
rect 894 42439 900 42442
rect 1548 42442 1584 42448
rect 1548 42439 1554 42442
rect 156 42402 162 42405
rect 126 42396 162 42402
rect 810 42402 816 42405
rect 810 42396 1584 42402
rect 126 42362 138 42396
rect 1572 42362 1584 42396
rect 126 42356 162 42362
rect 156 42353 162 42356
rect 810 42356 1584 42362
rect 810 42353 816 42356
rect 894 42316 900 42319
rect 126 42310 900 42316
rect 1548 42316 1554 42319
rect 1548 42310 1584 42316
rect 126 42276 138 42310
rect 1572 42276 1584 42310
rect 126 42270 900 42276
rect 894 42267 900 42270
rect 1548 42270 1584 42276
rect 1548 42267 1554 42270
rect 156 42230 162 42233
rect 126 42224 162 42230
rect 810 42230 816 42233
rect 810 42224 1584 42230
rect 126 42190 138 42224
rect 1572 42190 1584 42224
rect 126 42184 162 42190
rect 156 42181 162 42184
rect 810 42184 1584 42190
rect 810 42181 816 42184
rect 894 42144 900 42147
rect 126 42138 900 42144
rect 1548 42144 1554 42147
rect 1548 42138 1584 42144
rect 126 42104 138 42138
rect 1572 42104 1584 42138
rect 126 42098 900 42104
rect 894 42095 900 42098
rect 1548 42098 1584 42104
rect 1548 42095 1554 42098
rect 156 42058 162 42061
rect 126 42052 162 42058
rect 810 42058 816 42061
rect 810 42052 1584 42058
rect 126 42018 138 42052
rect 1572 42018 1584 42052
rect 126 42012 162 42018
rect 156 42009 162 42012
rect 810 42012 1584 42018
rect 810 42009 816 42012
rect 894 41972 900 41975
rect 126 41966 900 41972
rect 1548 41972 1554 41975
rect 1548 41966 1584 41972
rect 126 41932 138 41966
rect 1572 41932 1584 41966
rect 126 41926 900 41932
rect 894 41923 900 41926
rect 1548 41926 1584 41932
rect 1548 41923 1554 41926
rect 156 41886 162 41889
rect 126 41880 162 41886
rect 810 41886 816 41889
rect 810 41880 1584 41886
rect 126 41846 138 41880
rect 1572 41846 1584 41880
rect 126 41840 162 41846
rect 156 41837 162 41840
rect 810 41840 1584 41846
rect 810 41837 816 41840
rect 894 41800 900 41803
rect 126 41794 900 41800
rect 1548 41800 1554 41803
rect 1548 41794 1584 41800
rect 126 41760 138 41794
rect 1572 41760 1584 41794
rect 126 41754 900 41760
rect 894 41751 900 41754
rect 1548 41754 1584 41760
rect 1548 41751 1554 41754
rect 156 41714 162 41717
rect 126 41708 162 41714
rect 810 41714 816 41717
rect 810 41708 1584 41714
rect 126 41674 138 41708
rect 1572 41674 1584 41708
rect 126 41668 162 41674
rect 156 41665 162 41668
rect 810 41668 1584 41674
rect 810 41665 816 41668
rect 894 41628 900 41631
rect 126 41622 900 41628
rect 1548 41628 1554 41631
rect 1548 41622 1584 41628
rect 126 41588 138 41622
rect 1572 41588 1584 41622
rect 126 41582 900 41588
rect 894 41579 900 41582
rect 1548 41582 1584 41588
rect 1548 41579 1554 41582
rect 156 41542 162 41545
rect 126 41536 162 41542
rect 810 41542 816 41545
rect 810 41536 1584 41542
rect 126 41502 138 41536
rect 1572 41502 1584 41536
rect 126 41496 162 41502
rect 156 41493 162 41496
rect 810 41496 1584 41502
rect 810 41493 816 41496
rect 894 41456 900 41459
rect 126 41450 900 41456
rect 1548 41456 1554 41459
rect 1548 41450 1584 41456
rect 126 41416 138 41450
rect 1572 41416 1584 41450
rect 126 41410 900 41416
rect 894 41407 900 41410
rect 1548 41410 1584 41416
rect 1548 41407 1554 41410
rect 156 41370 162 41373
rect 126 41364 162 41370
rect 810 41370 816 41373
rect 810 41364 1584 41370
rect 126 41330 138 41364
rect 1572 41330 1584 41364
rect 126 41324 162 41330
rect 156 41321 162 41324
rect 810 41324 1584 41330
rect 810 41321 816 41324
rect 894 41284 900 41287
rect 126 41278 900 41284
rect 1548 41284 1554 41287
rect 1548 41278 1584 41284
rect 126 41244 138 41278
rect 1572 41244 1584 41278
rect 126 41238 900 41244
rect 894 41235 900 41238
rect 1548 41238 1584 41244
rect 1548 41235 1554 41238
rect 156 41198 162 41201
rect 126 41192 162 41198
rect 810 41198 816 41201
rect 810 41192 1584 41198
rect 126 41158 138 41192
rect 1572 41158 1584 41192
rect 126 41152 162 41158
rect 156 41149 162 41152
rect 810 41152 1584 41158
rect 810 41149 816 41152
rect 894 41112 900 41115
rect 126 41106 900 41112
rect 1548 41112 1554 41115
rect 1548 41106 1584 41112
rect 126 41072 138 41106
rect 1572 41072 1584 41106
rect 126 41066 900 41072
rect 894 41063 900 41066
rect 1548 41066 1584 41072
rect 1548 41063 1554 41066
rect 156 41026 162 41029
rect 126 41020 162 41026
rect 810 41026 816 41029
rect 810 41020 1584 41026
rect 126 40986 138 41020
rect 1572 40986 1584 41020
rect 126 40980 162 40986
rect 156 40977 162 40980
rect 810 40980 1584 40986
rect 810 40977 816 40980
rect 894 40940 900 40943
rect 126 40934 900 40940
rect 1548 40940 1554 40943
rect 1548 40934 1584 40940
rect 126 40900 138 40934
rect 1572 40900 1584 40934
rect 126 40894 900 40900
rect 894 40891 900 40894
rect 1548 40894 1584 40900
rect 1548 40891 1554 40894
rect 156 40854 162 40857
rect 126 40848 162 40854
rect 810 40854 816 40857
rect 810 40848 1584 40854
rect 126 40814 138 40848
rect 1572 40814 1584 40848
rect 126 40808 162 40814
rect 156 40805 162 40808
rect 810 40808 1584 40814
rect 810 40805 816 40808
rect 894 40768 900 40771
rect 126 40762 900 40768
rect 1548 40768 1554 40771
rect 1548 40762 1584 40768
rect 126 40728 138 40762
rect 1572 40728 1584 40762
rect 126 40722 900 40728
rect 894 40719 900 40722
rect 1548 40722 1584 40728
rect 1548 40719 1554 40722
rect 156 40682 162 40685
rect 126 40676 162 40682
rect 810 40682 816 40685
rect 810 40676 1584 40682
rect 126 40642 138 40676
rect 1572 40642 1584 40676
rect 126 40636 162 40642
rect 156 40633 162 40636
rect 810 40636 1584 40642
rect 810 40633 816 40636
rect 894 40596 900 40599
rect 126 40590 900 40596
rect 1548 40596 1554 40599
rect 1548 40590 1584 40596
rect 126 40556 138 40590
rect 1572 40556 1584 40590
rect 126 40550 900 40556
rect 894 40547 900 40550
rect 1548 40550 1584 40556
rect 1548 40547 1554 40550
rect 156 40510 162 40513
rect 126 40504 162 40510
rect 810 40510 816 40513
rect 810 40504 1584 40510
rect 126 40470 138 40504
rect 1572 40470 1584 40504
rect 126 40464 162 40470
rect 156 40461 162 40464
rect 810 40464 1584 40470
rect 810 40461 816 40464
rect 894 40424 900 40427
rect 126 40418 900 40424
rect 1548 40424 1554 40427
rect 1548 40418 1584 40424
rect 126 40384 138 40418
rect 1572 40384 1584 40418
rect 126 40378 900 40384
rect 894 40375 900 40378
rect 1548 40378 1584 40384
rect 1548 40375 1554 40378
rect 156 40338 162 40341
rect 126 40332 162 40338
rect 810 40338 816 40341
rect 810 40332 1584 40338
rect 126 40298 138 40332
rect 1572 40298 1584 40332
rect 126 40292 162 40298
rect 156 40289 162 40292
rect 810 40292 1584 40298
rect 810 40289 816 40292
rect 894 40252 900 40255
rect 126 40246 900 40252
rect 1548 40252 1554 40255
rect 1548 40246 1584 40252
rect 126 40212 138 40246
rect 1572 40212 1584 40246
rect 126 40206 900 40212
rect 894 40203 900 40206
rect 1548 40206 1584 40212
rect 1548 40203 1554 40206
rect 156 40166 162 40169
rect 126 40160 162 40166
rect 810 40166 816 40169
rect 810 40160 1584 40166
rect 126 40126 138 40160
rect 1572 40126 1584 40160
rect 126 40120 162 40126
rect 156 40117 162 40120
rect 810 40120 1584 40126
rect 810 40117 816 40120
rect 894 40080 900 40083
rect 126 40074 900 40080
rect 1548 40080 1554 40083
rect 1548 40074 1584 40080
rect 126 40040 138 40074
rect 1572 40040 1584 40074
rect 126 40034 900 40040
rect 894 40031 900 40034
rect 1548 40034 1584 40040
rect 1548 40031 1554 40034
rect 156 39994 162 39997
rect 126 39988 162 39994
rect 810 39994 816 39997
rect 810 39988 1584 39994
rect 126 39954 138 39988
rect 1572 39954 1584 39988
rect 126 39948 162 39954
rect 156 39945 162 39948
rect 810 39948 1584 39954
rect 810 39945 816 39948
rect 894 39908 900 39911
rect 126 39902 900 39908
rect 1548 39908 1554 39911
rect 1548 39902 1584 39908
rect 126 39868 138 39902
rect 1572 39868 1584 39902
rect 126 39862 900 39868
rect 894 39859 900 39862
rect 1548 39862 1584 39868
rect 1548 39859 1554 39862
rect 156 39822 162 39825
rect 126 39816 162 39822
rect 810 39822 816 39825
rect 810 39816 1584 39822
rect 126 39782 138 39816
rect 1572 39782 1584 39816
rect 126 39776 162 39782
rect 156 39773 162 39776
rect 810 39776 1584 39782
rect 810 39773 816 39776
rect 894 39736 900 39739
rect 126 39730 900 39736
rect 1548 39736 1554 39739
rect 1548 39730 1584 39736
rect 126 39696 138 39730
rect 1572 39696 1584 39730
rect 126 39690 900 39696
rect 894 39687 900 39690
rect 1548 39690 1584 39696
rect 1548 39687 1554 39690
rect 156 39650 162 39653
rect 126 39644 162 39650
rect 810 39650 816 39653
rect 810 39644 1584 39650
rect 126 39610 138 39644
rect 1572 39610 1584 39644
rect 126 39604 162 39610
rect 156 39601 162 39604
rect 810 39604 1584 39610
rect 810 39601 816 39604
rect 894 39564 900 39567
rect 126 39558 900 39564
rect 1548 39564 1554 39567
rect 1548 39558 1584 39564
rect 126 39524 138 39558
rect 1572 39524 1584 39558
rect 126 39518 900 39524
rect 894 39515 900 39518
rect 1548 39518 1584 39524
rect 1548 39515 1554 39518
rect 156 39478 162 39481
rect 126 39472 162 39478
rect 810 39478 816 39481
rect 810 39472 1584 39478
rect 126 39438 138 39472
rect 1572 39438 1584 39472
rect 126 39432 162 39438
rect 156 39429 162 39432
rect 810 39432 1584 39438
rect 810 39429 816 39432
rect 894 39392 900 39395
rect 126 39386 900 39392
rect 1548 39392 1554 39395
rect 1548 39386 1584 39392
rect 126 39352 138 39386
rect 1572 39352 1584 39386
rect 126 39346 900 39352
rect 894 39343 900 39346
rect 1548 39346 1584 39352
rect 1548 39343 1554 39346
rect 156 39306 162 39309
rect 126 39300 162 39306
rect 810 39306 816 39309
rect 810 39300 1584 39306
rect 126 39266 138 39300
rect 1572 39266 1584 39300
rect 126 39260 162 39266
rect 156 39257 162 39260
rect 810 39260 1584 39266
rect 810 39257 816 39260
rect 894 39220 900 39223
rect 126 39214 900 39220
rect 1548 39220 1554 39223
rect 1548 39214 1584 39220
rect 126 39180 138 39214
rect 1572 39180 1584 39214
rect 126 39174 900 39180
rect 894 39171 900 39174
rect 1548 39174 1584 39180
rect 1548 39171 1554 39174
rect 156 39134 162 39137
rect 126 39128 162 39134
rect 810 39134 816 39137
rect 810 39128 1584 39134
rect 126 39094 138 39128
rect 1572 39094 1584 39128
rect 126 39088 162 39094
rect 156 39085 162 39088
rect 810 39088 1584 39094
rect 810 39085 816 39088
rect 894 39048 900 39051
rect 126 39042 900 39048
rect 1548 39048 1554 39051
rect 1548 39042 1584 39048
rect 126 39008 138 39042
rect 1572 39008 1584 39042
rect 126 39002 900 39008
rect 894 38999 900 39002
rect 1548 39002 1584 39008
rect 1548 38999 1554 39002
rect 156 38962 162 38965
rect 126 38956 162 38962
rect 810 38962 816 38965
rect 810 38956 1584 38962
rect 126 38922 138 38956
rect 1572 38922 1584 38956
rect 126 38916 162 38922
rect 156 38913 162 38916
rect 810 38916 1584 38922
rect 810 38913 816 38916
rect 894 38876 900 38879
rect 126 38870 900 38876
rect 1548 38876 1554 38879
rect 1548 38870 1584 38876
rect 126 38836 138 38870
rect 1572 38836 1584 38870
rect 126 38830 900 38836
rect 894 38827 900 38830
rect 1548 38830 1584 38836
rect 1548 38827 1554 38830
rect 156 38790 162 38793
rect 126 38784 162 38790
rect 810 38790 816 38793
rect 810 38784 1584 38790
rect 126 38750 138 38784
rect 1572 38750 1584 38784
rect 126 38744 162 38750
rect 156 38741 162 38744
rect 810 38744 1584 38750
rect 810 38741 816 38744
rect 894 38704 900 38707
rect 126 38698 900 38704
rect 1548 38704 1554 38707
rect 1548 38698 1584 38704
rect 126 38664 138 38698
rect 1572 38664 1584 38698
rect 126 38658 900 38664
rect 894 38655 900 38658
rect 1548 38658 1584 38664
rect 1548 38655 1554 38658
rect 156 38618 162 38621
rect 126 38612 162 38618
rect 810 38618 816 38621
rect 810 38612 1584 38618
rect 126 38578 138 38612
rect 1572 38578 1584 38612
rect 126 38572 162 38578
rect 156 38569 162 38572
rect 810 38572 1584 38578
rect 810 38569 816 38572
rect 894 38532 900 38535
rect 126 38526 900 38532
rect 1548 38532 1554 38535
rect 1548 38526 1584 38532
rect 126 38492 138 38526
rect 1572 38492 1584 38526
rect 126 38486 900 38492
rect 894 38483 900 38486
rect 1548 38486 1584 38492
rect 1548 38483 1554 38486
rect 156 38446 162 38449
rect 126 38440 162 38446
rect 810 38446 816 38449
rect 810 38440 1584 38446
rect 126 38406 138 38440
rect 1572 38406 1584 38440
rect 126 38400 162 38406
rect 156 38397 162 38400
rect 810 38400 1584 38406
rect 810 38397 816 38400
rect 894 38360 900 38363
rect 126 38354 900 38360
rect 1548 38360 1554 38363
rect 1548 38354 1584 38360
rect 126 38320 138 38354
rect 1572 38320 1584 38354
rect 126 38314 900 38320
rect 894 38311 900 38314
rect 1548 38314 1584 38320
rect 1548 38311 1554 38314
rect 156 38274 162 38277
rect 126 38268 162 38274
rect 810 38274 816 38277
rect 810 38268 1584 38274
rect 126 38234 138 38268
rect 1572 38234 1584 38268
rect 126 38228 162 38234
rect 156 38225 162 38228
rect 810 38228 1584 38234
rect 810 38225 816 38228
rect 894 38188 900 38191
rect 126 38182 900 38188
rect 1548 38188 1554 38191
rect 1548 38182 1584 38188
rect 126 38148 138 38182
rect 1572 38148 1584 38182
rect 126 38142 900 38148
rect 894 38139 900 38142
rect 1548 38142 1584 38148
rect 1548 38139 1554 38142
rect 156 38102 162 38105
rect 126 38096 162 38102
rect 810 38102 816 38105
rect 810 38096 1584 38102
rect 126 38062 138 38096
rect 1572 38062 1584 38096
rect 126 38056 162 38062
rect 156 38053 162 38056
rect 810 38056 1584 38062
rect 810 38053 816 38056
rect 894 38016 900 38019
rect 126 38010 900 38016
rect 1548 38016 1554 38019
rect 1548 38010 1584 38016
rect 126 37976 138 38010
rect 1572 37976 1584 38010
rect 126 37970 900 37976
rect 894 37967 900 37970
rect 1548 37970 1584 37976
rect 1548 37967 1554 37970
rect 156 37930 162 37933
rect 126 37924 162 37930
rect 810 37930 816 37933
rect 810 37924 1584 37930
rect 126 37890 138 37924
rect 1572 37890 1584 37924
rect 126 37884 162 37890
rect 156 37881 162 37884
rect 810 37884 1584 37890
rect 810 37881 816 37884
rect 894 37844 900 37847
rect 126 37838 900 37844
rect 1548 37844 1554 37847
rect 1548 37838 1584 37844
rect 126 37804 138 37838
rect 1572 37804 1584 37838
rect 126 37798 900 37804
rect 894 37795 900 37798
rect 1548 37798 1584 37804
rect 1548 37795 1554 37798
rect 156 37758 162 37761
rect 126 37752 162 37758
rect 810 37758 816 37761
rect 810 37752 1584 37758
rect 126 37718 138 37752
rect 1572 37718 1584 37752
rect 126 37712 162 37718
rect 156 37709 162 37712
rect 810 37712 1584 37718
rect 810 37709 816 37712
rect 894 37672 900 37675
rect 126 37666 900 37672
rect 1548 37672 1554 37675
rect 1548 37666 1584 37672
rect 126 37632 138 37666
rect 1572 37632 1584 37666
rect 126 37626 900 37632
rect 894 37623 900 37626
rect 1548 37626 1584 37632
rect 1548 37623 1554 37626
rect 156 37586 162 37589
rect 126 37580 162 37586
rect 810 37586 816 37589
rect 810 37580 1584 37586
rect 126 37546 138 37580
rect 1572 37546 1584 37580
rect 126 37540 162 37546
rect 156 37537 162 37540
rect 810 37540 1584 37546
rect 810 37537 816 37540
rect 894 37500 900 37503
rect 126 37494 900 37500
rect 1548 37500 1554 37503
rect 1548 37494 1584 37500
rect 126 37460 138 37494
rect 1572 37460 1584 37494
rect 126 37454 900 37460
rect 894 37451 900 37454
rect 1548 37454 1584 37460
rect 1548 37451 1554 37454
rect 156 37414 162 37417
rect 126 37408 162 37414
rect 810 37414 816 37417
rect 810 37408 1584 37414
rect 126 37374 138 37408
rect 1572 37374 1584 37408
rect 126 37368 162 37374
rect 156 37365 162 37368
rect 810 37368 1584 37374
rect 810 37365 816 37368
rect 894 37328 900 37331
rect 126 37322 900 37328
rect 1548 37328 1554 37331
rect 1548 37322 1584 37328
rect 126 37288 138 37322
rect 1572 37288 1584 37322
rect 126 37282 900 37288
rect 894 37279 900 37282
rect 1548 37282 1584 37288
rect 1548 37279 1554 37282
rect 156 37242 162 37245
rect 126 37236 162 37242
rect 810 37242 816 37245
rect 810 37236 1584 37242
rect 126 37202 138 37236
rect 1572 37202 1584 37236
rect 126 37196 162 37202
rect 156 37193 162 37196
rect 810 37196 1584 37202
rect 810 37193 816 37196
rect 894 37156 900 37159
rect 126 37150 900 37156
rect 1548 37156 1554 37159
rect 1548 37150 1584 37156
rect 126 37116 138 37150
rect 1572 37116 1584 37150
rect 126 37110 900 37116
rect 894 37107 900 37110
rect 1548 37110 1584 37116
rect 1548 37107 1554 37110
rect 156 37070 162 37073
rect 126 37064 162 37070
rect 810 37070 816 37073
rect 810 37064 1584 37070
rect 126 37030 138 37064
rect 1572 37030 1584 37064
rect 126 37024 162 37030
rect 156 37021 162 37024
rect 810 37024 1584 37030
rect 810 37021 816 37024
rect 894 36984 900 36987
rect 126 36978 900 36984
rect 1548 36984 1554 36987
rect 1548 36978 1584 36984
rect 126 36944 138 36978
rect 1572 36944 1584 36978
rect 126 36938 900 36944
rect 894 36935 900 36938
rect 1548 36938 1584 36944
rect 1548 36935 1554 36938
rect 156 36898 162 36901
rect 126 36892 162 36898
rect 810 36898 816 36901
rect 810 36892 1584 36898
rect 126 36858 138 36892
rect 1572 36858 1584 36892
rect 126 36852 162 36858
rect 156 36849 162 36852
rect 810 36852 1584 36858
rect 810 36849 816 36852
rect 894 36812 900 36815
rect 126 36806 900 36812
rect 1548 36812 1554 36815
rect 1548 36806 1584 36812
rect 126 36772 138 36806
rect 1572 36772 1584 36806
rect 126 36766 900 36772
rect 894 36763 900 36766
rect 1548 36766 1584 36772
rect 1548 36763 1554 36766
rect 156 36726 162 36729
rect 126 36720 162 36726
rect 810 36726 816 36729
rect 810 36720 1584 36726
rect 126 36686 138 36720
rect 1572 36686 1584 36720
rect 126 36680 162 36686
rect 156 36677 162 36680
rect 810 36680 1584 36686
rect 810 36677 816 36680
rect 894 36640 900 36643
rect 126 36634 900 36640
rect 1548 36640 1554 36643
rect 1548 36634 1584 36640
rect 126 36600 138 36634
rect 1572 36600 1584 36634
rect 126 36594 900 36600
rect 894 36591 900 36594
rect 1548 36594 1584 36600
rect 1548 36591 1554 36594
rect 156 36554 162 36557
rect 126 36548 162 36554
rect 810 36554 816 36557
rect 810 36548 1584 36554
rect 126 36514 138 36548
rect 1572 36514 1584 36548
rect 126 36508 162 36514
rect 156 36505 162 36508
rect 810 36508 1584 36514
rect 810 36505 816 36508
rect 894 36468 900 36471
rect 126 36462 900 36468
rect 1548 36468 1554 36471
rect 1548 36462 1584 36468
rect 126 36428 138 36462
rect 1572 36428 1584 36462
rect 126 36422 900 36428
rect 894 36419 900 36422
rect 1548 36422 1584 36428
rect 1548 36419 1554 36422
rect 156 36382 162 36385
rect 126 36376 162 36382
rect 810 36382 816 36385
rect 810 36376 1584 36382
rect 126 36342 138 36376
rect 1572 36342 1584 36376
rect 126 36336 162 36342
rect 156 36333 162 36336
rect 810 36336 1584 36342
rect 810 36333 816 36336
rect 894 36296 900 36299
rect 126 36290 900 36296
rect 1548 36296 1554 36299
rect 1548 36290 1584 36296
rect 126 36256 138 36290
rect 1572 36256 1584 36290
rect 126 36250 900 36256
rect 894 36247 900 36250
rect 1548 36250 1584 36256
rect 1548 36247 1554 36250
rect 156 36210 162 36213
rect 126 36204 162 36210
rect 810 36210 816 36213
rect 810 36204 1584 36210
rect 126 36170 138 36204
rect 1572 36170 1584 36204
rect 126 36164 162 36170
rect 156 36161 162 36164
rect 810 36164 1584 36170
rect 810 36161 816 36164
rect 894 36124 900 36127
rect 126 36118 900 36124
rect 1548 36124 1554 36127
rect 1548 36118 1584 36124
rect 126 36084 138 36118
rect 1572 36084 1584 36118
rect 126 36078 900 36084
rect 894 36075 900 36078
rect 1548 36078 1584 36084
rect 1548 36075 1554 36078
rect 156 36038 162 36041
rect 126 36032 162 36038
rect 810 36038 816 36041
rect 810 36032 1584 36038
rect 126 35998 138 36032
rect 1572 35998 1584 36032
rect 126 35992 162 35998
rect 156 35989 162 35992
rect 810 35992 1584 35998
rect 810 35989 816 35992
rect 894 35952 900 35955
rect 126 35946 900 35952
rect 1548 35952 1554 35955
rect 1548 35946 1584 35952
rect 126 35912 138 35946
rect 1572 35912 1584 35946
rect 126 35906 900 35912
rect 894 35903 900 35906
rect 1548 35906 1584 35912
rect 1548 35903 1554 35906
rect 156 35866 162 35869
rect 126 35860 162 35866
rect 810 35866 816 35869
rect 810 35860 1584 35866
rect 126 35826 138 35860
rect 1572 35826 1584 35860
rect 126 35820 162 35826
rect 156 35817 162 35820
rect 810 35820 1584 35826
rect 810 35817 816 35820
rect 894 35780 900 35783
rect 126 35774 900 35780
rect 1548 35780 1554 35783
rect 1548 35774 1584 35780
rect 126 35740 138 35774
rect 1572 35740 1584 35774
rect 126 35734 900 35740
rect 894 35731 900 35734
rect 1548 35734 1584 35740
rect 1548 35731 1554 35734
rect 156 35694 162 35697
rect 126 35688 162 35694
rect 810 35694 816 35697
rect 810 35688 1584 35694
rect 126 35654 138 35688
rect 1572 35654 1584 35688
rect 126 35648 162 35654
rect 156 35645 162 35648
rect 810 35648 1584 35654
rect 810 35645 816 35648
rect 894 35608 900 35611
rect 126 35602 900 35608
rect 1548 35608 1554 35611
rect 1548 35602 1584 35608
rect 126 35568 138 35602
rect 1572 35568 1584 35602
rect 126 35562 900 35568
rect 894 35559 900 35562
rect 1548 35562 1584 35568
rect 1548 35559 1554 35562
rect 156 35522 162 35525
rect 126 35516 162 35522
rect 810 35522 816 35525
rect 810 35516 1584 35522
rect 126 35482 138 35516
rect 1572 35482 1584 35516
rect 126 35476 162 35482
rect 156 35473 162 35476
rect 810 35476 1584 35482
rect 810 35473 816 35476
rect 894 35436 900 35439
rect 126 35430 900 35436
rect 1548 35436 1554 35439
rect 1548 35430 1584 35436
rect 126 35396 138 35430
rect 1572 35396 1584 35430
rect 126 35390 900 35396
rect 894 35387 900 35390
rect 1548 35390 1584 35396
rect 1548 35387 1554 35390
rect 156 35350 162 35353
rect 126 35344 162 35350
rect 810 35350 816 35353
rect 810 35344 1584 35350
rect 126 35310 138 35344
rect 1572 35310 1584 35344
rect 126 35304 162 35310
rect 156 35301 162 35304
rect 810 35304 1584 35310
rect 810 35301 816 35304
rect 894 35264 900 35267
rect 126 35258 900 35264
rect 1548 35264 1554 35267
rect 1548 35258 1584 35264
rect 126 35224 138 35258
rect 1572 35224 1584 35258
rect 126 35218 900 35224
rect 894 35215 900 35218
rect 1548 35218 1584 35224
rect 1548 35215 1554 35218
rect 156 35178 162 35181
rect 126 35172 162 35178
rect 810 35178 816 35181
rect 810 35172 1584 35178
rect 126 35138 138 35172
rect 1572 35138 1584 35172
rect 126 35132 162 35138
rect 156 35129 162 35132
rect 810 35132 1584 35138
rect 810 35129 816 35132
rect 894 35092 900 35095
rect 126 35086 900 35092
rect 1548 35092 1554 35095
rect 1548 35086 1584 35092
rect 126 35052 138 35086
rect 1572 35052 1584 35086
rect 126 35046 900 35052
rect 894 35043 900 35046
rect 1548 35046 1584 35052
rect 1548 35043 1554 35046
rect 156 35006 162 35009
rect 126 35000 162 35006
rect 810 35006 816 35009
rect 810 35000 1584 35006
rect 126 34966 138 35000
rect 1572 34966 1584 35000
rect 126 34960 162 34966
rect 156 34957 162 34960
rect 810 34960 1584 34966
rect 810 34957 816 34960
rect 894 34920 900 34923
rect 126 34914 900 34920
rect 1548 34920 1554 34923
rect 1548 34914 1584 34920
rect 126 34880 138 34914
rect 1572 34880 1584 34914
rect 126 34874 900 34880
rect 894 34871 900 34874
rect 1548 34874 1584 34880
rect 1548 34871 1554 34874
rect 156 34834 162 34837
rect 126 34828 162 34834
rect 810 34834 816 34837
rect 810 34828 1584 34834
rect 126 34794 138 34828
rect 1572 34794 1584 34828
rect 126 34788 162 34794
rect 156 34785 162 34788
rect 810 34788 1584 34794
rect 810 34785 816 34788
rect 894 34748 900 34751
rect 126 34742 900 34748
rect 1548 34748 1554 34751
rect 1548 34742 1584 34748
rect 126 34708 138 34742
rect 1572 34708 1584 34742
rect 126 34702 900 34708
rect 894 34699 900 34702
rect 1548 34702 1584 34708
rect 1548 34699 1554 34702
rect 156 34662 162 34665
rect 126 34656 162 34662
rect 810 34662 816 34665
rect 810 34656 1584 34662
rect 126 34622 138 34656
rect 1572 34622 1584 34656
rect 126 34616 162 34622
rect 156 34613 162 34616
rect 810 34616 1584 34622
rect 810 34613 816 34616
rect 894 34576 900 34579
rect 126 34570 900 34576
rect 1548 34576 1554 34579
rect 1548 34570 1584 34576
rect 126 34536 138 34570
rect 1572 34536 1584 34570
rect 126 34530 900 34536
rect 894 34527 900 34530
rect 1548 34530 1584 34536
rect 1548 34527 1554 34530
rect 156 34490 162 34493
rect 126 34484 162 34490
rect 810 34490 816 34493
rect 810 34484 1584 34490
rect 126 34450 138 34484
rect 1572 34450 1584 34484
rect 126 34444 162 34450
rect 156 34441 162 34444
rect 810 34444 1584 34450
rect 810 34441 816 34444
rect 894 34404 900 34407
rect 126 34398 900 34404
rect 1548 34404 1554 34407
rect 1548 34398 1584 34404
rect 126 34364 138 34398
rect 1572 34364 1584 34398
rect 126 34358 900 34364
rect 894 34355 900 34358
rect 1548 34358 1584 34364
rect 1548 34355 1554 34358
rect 156 34318 162 34321
rect 126 34312 162 34318
rect 810 34318 816 34321
rect 810 34312 1584 34318
rect 126 34278 138 34312
rect 1572 34278 1584 34312
rect 126 34272 162 34278
rect 156 34269 162 34272
rect 810 34272 1584 34278
rect 810 34269 816 34272
rect 894 34232 900 34235
rect 126 34226 900 34232
rect 1548 34232 1554 34235
rect 1548 34226 1584 34232
rect 126 34192 138 34226
rect 1572 34192 1584 34226
rect 126 34186 900 34192
rect 894 34183 900 34186
rect 1548 34186 1584 34192
rect 1548 34183 1554 34186
rect 156 34146 162 34149
rect 126 34140 162 34146
rect 810 34146 816 34149
rect 810 34140 1584 34146
rect 126 34106 138 34140
rect 1572 34106 1584 34140
rect 126 34100 162 34106
rect 156 34097 162 34100
rect 810 34100 1584 34106
rect 810 34097 816 34100
rect 894 34060 900 34063
rect 126 34054 900 34060
rect 1548 34060 1554 34063
rect 1548 34054 1584 34060
rect 126 34020 138 34054
rect 1572 34020 1584 34054
rect 126 34014 900 34020
rect 894 34011 900 34014
rect 1548 34014 1584 34020
rect 1548 34011 1554 34014
rect 156 33974 162 33977
rect 126 33968 162 33974
rect 810 33974 816 33977
rect 810 33968 1584 33974
rect 126 33934 138 33968
rect 1572 33934 1584 33968
rect 126 33928 162 33934
rect 156 33925 162 33928
rect 810 33928 1584 33934
rect 810 33925 816 33928
rect 894 33888 900 33891
rect 126 33882 900 33888
rect 1548 33888 1554 33891
rect 1548 33882 1584 33888
rect 126 33848 138 33882
rect 1572 33848 1584 33882
rect 126 33842 900 33848
rect 894 33839 900 33842
rect 1548 33842 1584 33848
rect 1548 33839 1554 33842
rect 156 33802 162 33805
rect 126 33796 162 33802
rect 810 33802 816 33805
rect 810 33796 1584 33802
rect 126 33762 138 33796
rect 1572 33762 1584 33796
rect 126 33756 162 33762
rect 156 33753 162 33756
rect 810 33756 1584 33762
rect 810 33753 816 33756
rect 894 33716 900 33719
rect 126 33710 900 33716
rect 1548 33716 1554 33719
rect 1548 33710 1584 33716
rect 126 33676 138 33710
rect 1572 33676 1584 33710
rect 126 33670 900 33676
rect 894 33667 900 33670
rect 1548 33670 1584 33676
rect 1548 33667 1554 33670
rect 156 33630 162 33633
rect 126 33624 162 33630
rect 810 33630 816 33633
rect 810 33624 1584 33630
rect 126 33590 138 33624
rect 1572 33590 1584 33624
rect 126 33584 162 33590
rect 156 33581 162 33584
rect 810 33584 1584 33590
rect 810 33581 816 33584
rect 894 33544 900 33547
rect 126 33538 900 33544
rect 1548 33544 1554 33547
rect 1548 33538 1584 33544
rect 126 33504 138 33538
rect 1572 33504 1584 33538
rect 126 33498 900 33504
rect 894 33495 900 33498
rect 1548 33498 1584 33504
rect 1548 33495 1554 33498
rect 156 33458 162 33461
rect 126 33452 162 33458
rect 810 33458 816 33461
rect 810 33452 1584 33458
rect 126 33418 138 33452
rect 1572 33418 1584 33452
rect 126 33412 162 33418
rect 156 33409 162 33412
rect 810 33412 1584 33418
rect 810 33409 816 33412
rect 894 33372 900 33375
rect 126 33366 900 33372
rect 1548 33372 1554 33375
rect 1548 33366 1584 33372
rect 126 33332 138 33366
rect 1572 33332 1584 33366
rect 126 33326 900 33332
rect 894 33323 900 33326
rect 1548 33326 1584 33332
rect 1548 33323 1554 33326
rect 156 33286 162 33289
rect 126 33280 162 33286
rect 810 33286 816 33289
rect 810 33280 1584 33286
rect 126 33246 138 33280
rect 1572 33246 1584 33280
rect 126 33240 162 33246
rect 156 33237 162 33240
rect 810 33240 1584 33246
rect 810 33237 816 33240
rect 894 33200 900 33203
rect 126 33194 900 33200
rect 1548 33200 1554 33203
rect 1548 33194 1584 33200
rect 126 33160 138 33194
rect 1572 33160 1584 33194
rect 126 33154 900 33160
rect 894 33151 900 33154
rect 1548 33154 1584 33160
rect 1548 33151 1554 33154
rect 156 33114 162 33117
rect 126 33108 162 33114
rect 810 33114 816 33117
rect 810 33108 1584 33114
rect 126 33074 138 33108
rect 1572 33074 1584 33108
rect 126 33068 162 33074
rect 156 33065 162 33068
rect 810 33068 1584 33074
rect 810 33065 816 33068
rect 894 33028 900 33031
rect 126 33022 900 33028
rect 1548 33028 1554 33031
rect 1548 33022 1584 33028
rect 126 32988 138 33022
rect 1572 32988 1584 33022
rect 126 32982 900 32988
rect 894 32979 900 32982
rect 1548 32982 1584 32988
rect 1548 32979 1554 32982
rect 156 32942 162 32945
rect 126 32936 162 32942
rect 810 32942 816 32945
rect 810 32936 1584 32942
rect 126 32902 138 32936
rect 1572 32902 1584 32936
rect 126 32896 162 32902
rect 156 32893 162 32896
rect 810 32896 1584 32902
rect 810 32893 816 32896
rect 894 32856 900 32859
rect 126 32850 900 32856
rect 1548 32856 1554 32859
rect 1548 32850 1584 32856
rect 126 32816 138 32850
rect 1572 32816 1584 32850
rect 126 32810 900 32816
rect 894 32807 900 32810
rect 1548 32810 1584 32816
rect 1548 32807 1554 32810
rect 156 32770 162 32773
rect 126 32764 162 32770
rect 810 32770 816 32773
rect 810 32764 1584 32770
rect 126 32730 138 32764
rect 1572 32730 1584 32764
rect 126 32724 162 32730
rect 156 32721 162 32724
rect 810 32724 1584 32730
rect 810 32721 816 32724
rect 894 32684 900 32687
rect 126 32678 900 32684
rect 1548 32684 1554 32687
rect 1548 32678 1584 32684
rect 126 32644 138 32678
rect 1572 32644 1584 32678
rect 126 32638 900 32644
rect 894 32635 900 32638
rect 1548 32638 1584 32644
rect 1548 32635 1554 32638
rect 156 32598 162 32601
rect 126 32592 162 32598
rect 810 32598 816 32601
rect 810 32592 1584 32598
rect 126 32558 138 32592
rect 1572 32558 1584 32592
rect 126 32552 162 32558
rect 156 32549 162 32552
rect 810 32552 1584 32558
rect 810 32549 816 32552
rect 894 32512 900 32515
rect 126 32506 900 32512
rect 1548 32512 1554 32515
rect 1548 32506 1584 32512
rect 126 32472 138 32506
rect 1572 32472 1584 32506
rect 126 32466 900 32472
rect 894 32463 900 32466
rect 1548 32466 1584 32472
rect 1548 32463 1554 32466
rect 156 32426 162 32429
rect 126 32420 162 32426
rect 810 32426 816 32429
rect 810 32420 1584 32426
rect 126 32386 138 32420
rect 1572 32386 1584 32420
rect 126 32380 162 32386
rect 156 32377 162 32380
rect 810 32380 1584 32386
rect 810 32377 816 32380
rect 894 32340 900 32343
rect 126 32334 900 32340
rect 1548 32340 1554 32343
rect 1548 32334 1584 32340
rect 126 32300 138 32334
rect 1572 32300 1584 32334
rect 126 32294 900 32300
rect 894 32291 900 32294
rect 1548 32294 1584 32300
rect 1548 32291 1554 32294
rect 156 32254 162 32257
rect 126 32248 162 32254
rect 810 32254 816 32257
rect 810 32248 1584 32254
rect 126 32214 138 32248
rect 1572 32214 1584 32248
rect 126 32208 162 32214
rect 156 32205 162 32208
rect 810 32208 1584 32214
rect 810 32205 816 32208
rect 894 32168 900 32171
rect 126 32162 900 32168
rect 1548 32168 1554 32171
rect 1548 32162 1584 32168
rect 126 32128 138 32162
rect 1572 32128 1584 32162
rect 126 32122 900 32128
rect 894 32119 900 32122
rect 1548 32122 1584 32128
rect 1548 32119 1554 32122
rect 156 32082 162 32085
rect 126 32076 162 32082
rect 810 32082 816 32085
rect 810 32076 1584 32082
rect 126 32042 138 32076
rect 1572 32042 1584 32076
rect 126 32036 162 32042
rect 156 32033 162 32036
rect 810 32036 1584 32042
rect 810 32033 816 32036
rect 894 31996 900 31999
rect 126 31990 900 31996
rect 1548 31996 1554 31999
rect 1548 31990 1584 31996
rect 126 31956 138 31990
rect 1572 31956 1584 31990
rect 126 31950 900 31956
rect 894 31947 900 31950
rect 1548 31950 1584 31956
rect 1548 31947 1554 31950
rect 156 31910 162 31913
rect 126 31904 162 31910
rect 810 31910 816 31913
rect 810 31904 1584 31910
rect 126 31870 138 31904
rect 1572 31870 1584 31904
rect 126 31864 162 31870
rect 156 31861 162 31864
rect 810 31864 1584 31870
rect 810 31861 816 31864
rect 894 31824 900 31827
rect 126 31818 900 31824
rect 1548 31824 1554 31827
rect 1548 31818 1584 31824
rect 126 31784 138 31818
rect 1572 31784 1584 31818
rect 126 31778 900 31784
rect 894 31775 900 31778
rect 1548 31778 1584 31784
rect 1548 31775 1554 31778
rect 156 31738 162 31741
rect 126 31732 162 31738
rect 810 31738 816 31741
rect 810 31732 1584 31738
rect 126 31698 138 31732
rect 1572 31698 1584 31732
rect 126 31692 162 31698
rect 156 31689 162 31692
rect 810 31692 1584 31698
rect 810 31689 816 31692
rect 894 31652 900 31655
rect 126 31646 900 31652
rect 1548 31652 1554 31655
rect 1548 31646 1584 31652
rect 126 31612 138 31646
rect 1572 31612 1584 31646
rect 126 31606 900 31612
rect 894 31603 900 31606
rect 1548 31606 1584 31612
rect 1548 31603 1554 31606
rect 156 31566 162 31569
rect 126 31560 162 31566
rect 810 31566 816 31569
rect 810 31560 1584 31566
rect 126 31526 138 31560
rect 1572 31526 1584 31560
rect 126 31520 162 31526
rect 156 31517 162 31520
rect 810 31520 1584 31526
rect 810 31517 816 31520
rect 894 31480 900 31483
rect 126 31474 900 31480
rect 1548 31480 1554 31483
rect 1548 31474 1584 31480
rect 126 31440 138 31474
rect 1572 31440 1584 31474
rect 126 31434 900 31440
rect 894 31431 900 31434
rect 1548 31434 1584 31440
rect 1548 31431 1554 31434
rect 156 31394 162 31397
rect 126 31388 162 31394
rect 810 31394 816 31397
rect 810 31388 1584 31394
rect 126 31354 138 31388
rect 1572 31354 1584 31388
rect 126 31348 162 31354
rect 156 31345 162 31348
rect 810 31348 1584 31354
rect 810 31345 816 31348
rect 894 31308 900 31311
rect 126 31302 900 31308
rect 1548 31308 1554 31311
rect 1548 31302 1584 31308
rect 126 31268 138 31302
rect 1572 31268 1584 31302
rect 126 31262 900 31268
rect 894 31259 900 31262
rect 1548 31262 1584 31268
rect 1548 31259 1554 31262
rect 156 31222 162 31225
rect 126 31216 162 31222
rect 810 31222 816 31225
rect 810 31216 1584 31222
rect 126 31182 138 31216
rect 1572 31182 1584 31216
rect 126 31176 162 31182
rect 156 31173 162 31176
rect 810 31176 1584 31182
rect 810 31173 816 31176
rect 894 31136 900 31139
rect 126 31130 900 31136
rect 1548 31136 1554 31139
rect 1548 31130 1584 31136
rect 126 31096 138 31130
rect 1572 31096 1584 31130
rect 126 31090 900 31096
rect 894 31087 900 31090
rect 1548 31090 1584 31096
rect 1548 31087 1554 31090
rect 156 31050 162 31053
rect 126 31044 162 31050
rect 810 31050 816 31053
rect 810 31044 1584 31050
rect 126 31010 138 31044
rect 1572 31010 1584 31044
rect 126 31004 162 31010
rect 156 31001 162 31004
rect 810 31004 1584 31010
rect 810 31001 816 31004
rect 894 30964 900 30967
rect 126 30958 900 30964
rect 1548 30964 1554 30967
rect 1548 30958 1584 30964
rect 126 30924 138 30958
rect 1572 30924 1584 30958
rect 126 30918 900 30924
rect 894 30915 900 30918
rect 1548 30918 1584 30924
rect 1548 30915 1554 30918
rect 156 30878 162 30881
rect 126 30872 162 30878
rect 810 30878 816 30881
rect 810 30872 1584 30878
rect 126 30838 138 30872
rect 1572 30838 1584 30872
rect 126 30832 162 30838
rect 156 30829 162 30832
rect 810 30832 1584 30838
rect 810 30829 816 30832
rect 894 30792 900 30795
rect 126 30786 900 30792
rect 1548 30792 1554 30795
rect 1548 30786 1584 30792
rect 126 30752 138 30786
rect 1572 30752 1584 30786
rect 126 30746 900 30752
rect 894 30743 900 30746
rect 1548 30746 1584 30752
rect 1548 30743 1554 30746
rect 156 30706 162 30709
rect 126 30700 162 30706
rect 810 30706 816 30709
rect 810 30700 1584 30706
rect 126 30666 138 30700
rect 1572 30666 1584 30700
rect 126 30660 162 30666
rect 156 30657 162 30660
rect 810 30660 1584 30666
rect 810 30657 816 30660
rect 894 30620 900 30623
rect 126 30614 900 30620
rect 1548 30620 1554 30623
rect 1548 30614 1584 30620
rect 126 30580 138 30614
rect 1572 30580 1584 30614
rect 126 30574 900 30580
rect 894 30571 900 30574
rect 1548 30574 1584 30580
rect 1548 30571 1554 30574
rect 156 30534 162 30537
rect 126 30528 162 30534
rect 810 30534 816 30537
rect 810 30528 1584 30534
rect 126 30494 138 30528
rect 1572 30494 1584 30528
rect 126 30488 162 30494
rect 156 30485 162 30488
rect 810 30488 1584 30494
rect 810 30485 816 30488
rect 894 30448 900 30451
rect 126 30442 900 30448
rect 1548 30448 1554 30451
rect 1548 30442 1584 30448
rect 126 30408 138 30442
rect 1572 30408 1584 30442
rect 126 30402 900 30408
rect 894 30399 900 30402
rect 1548 30402 1584 30408
rect 1548 30399 1554 30402
rect 156 30362 162 30365
rect 126 30356 162 30362
rect 810 30362 816 30365
rect 810 30356 1584 30362
rect 126 30322 138 30356
rect 1572 30322 1584 30356
rect 126 30316 162 30322
rect 156 30313 162 30316
rect 810 30316 1584 30322
rect 810 30313 816 30316
rect 894 30276 900 30279
rect 126 30270 900 30276
rect 1548 30276 1554 30279
rect 1548 30270 1584 30276
rect 126 30236 138 30270
rect 1572 30236 1584 30270
rect 126 30230 900 30236
rect 894 30227 900 30230
rect 1548 30230 1584 30236
rect 1548 30227 1554 30230
rect 156 30190 162 30193
rect 126 30184 162 30190
rect 810 30190 816 30193
rect 810 30184 1584 30190
rect 126 30150 138 30184
rect 1572 30150 1584 30184
rect 126 30144 162 30150
rect 156 30141 162 30144
rect 810 30144 1584 30150
rect 810 30141 816 30144
rect 894 30104 900 30107
rect 126 30098 900 30104
rect 1548 30104 1554 30107
rect 1548 30098 1584 30104
rect 126 30064 138 30098
rect 1572 30064 1584 30098
rect 126 30058 900 30064
rect 894 30055 900 30058
rect 1548 30058 1584 30064
rect 1548 30055 1554 30058
rect 156 30018 162 30021
rect 126 30012 162 30018
rect 810 30018 816 30021
rect 810 30012 1584 30018
rect 126 29978 138 30012
rect 1572 29978 1584 30012
rect 126 29972 162 29978
rect 156 29969 162 29972
rect 810 29972 1584 29978
rect 810 29969 816 29972
rect 894 29932 900 29935
rect 126 29926 900 29932
rect 1548 29932 1554 29935
rect 1548 29926 1584 29932
rect 126 29892 138 29926
rect 1572 29892 1584 29926
rect 126 29886 900 29892
rect 894 29883 900 29886
rect 1548 29886 1584 29892
rect 1548 29883 1554 29886
rect 156 29846 162 29849
rect 126 29840 162 29846
rect 810 29846 816 29849
rect 810 29840 1584 29846
rect 126 29806 138 29840
rect 1572 29806 1584 29840
rect 126 29800 162 29806
rect 156 29797 162 29800
rect 810 29800 1584 29806
rect 810 29797 816 29800
rect 894 29760 900 29763
rect 126 29754 900 29760
rect 1548 29760 1554 29763
rect 1548 29754 1584 29760
rect 126 29720 138 29754
rect 1572 29720 1584 29754
rect 126 29714 900 29720
rect 894 29711 900 29714
rect 1548 29714 1584 29720
rect 1548 29711 1554 29714
rect 156 29674 162 29677
rect 126 29668 162 29674
rect 810 29674 816 29677
rect 810 29668 1584 29674
rect 126 29634 138 29668
rect 1572 29634 1584 29668
rect 126 29628 162 29634
rect 156 29625 162 29628
rect 810 29628 1584 29634
rect 810 29625 816 29628
rect 894 29588 900 29591
rect 126 29582 900 29588
rect 1548 29588 1554 29591
rect 1548 29582 1584 29588
rect 126 29548 138 29582
rect 1572 29548 1584 29582
rect 126 29542 900 29548
rect 894 29539 900 29542
rect 1548 29542 1584 29548
rect 1548 29539 1554 29542
rect 156 29502 162 29505
rect 126 29496 162 29502
rect 810 29502 816 29505
rect 810 29496 1584 29502
rect 126 29462 138 29496
rect 1572 29462 1584 29496
rect 126 29456 162 29462
rect 156 29453 162 29456
rect 810 29456 1584 29462
rect 810 29453 816 29456
rect 894 29416 900 29419
rect 126 29410 900 29416
rect 1548 29416 1554 29419
rect 1548 29410 1584 29416
rect 126 29376 138 29410
rect 1572 29376 1584 29410
rect 126 29370 900 29376
rect 894 29367 900 29370
rect 1548 29370 1584 29376
rect 1548 29367 1554 29370
rect 156 29330 162 29333
rect 126 29324 162 29330
rect 810 29330 816 29333
rect 810 29324 1584 29330
rect 126 29290 138 29324
rect 1572 29290 1584 29324
rect 126 29284 162 29290
rect 156 29281 162 29284
rect 810 29284 1584 29290
rect 810 29281 816 29284
rect 894 29244 900 29247
rect 126 29238 900 29244
rect 1548 29244 1554 29247
rect 1548 29238 1584 29244
rect 126 29204 138 29238
rect 1572 29204 1584 29238
rect 126 29198 900 29204
rect 894 29195 900 29198
rect 1548 29198 1584 29204
rect 1548 29195 1554 29198
rect 156 29158 162 29161
rect 126 29152 162 29158
rect 810 29158 816 29161
rect 810 29152 1584 29158
rect 126 29118 138 29152
rect 1572 29118 1584 29152
rect 126 29112 162 29118
rect 156 29109 162 29112
rect 810 29112 1584 29118
rect 810 29109 816 29112
rect 894 29072 900 29075
rect 126 29066 900 29072
rect 1548 29072 1554 29075
rect 1548 29066 1584 29072
rect 126 29032 138 29066
rect 1572 29032 1584 29066
rect 126 29026 900 29032
rect 894 29023 900 29026
rect 1548 29026 1584 29032
rect 1548 29023 1554 29026
rect 156 28986 162 28989
rect 126 28980 162 28986
rect 810 28986 816 28989
rect 810 28980 1584 28986
rect 126 28946 138 28980
rect 1572 28946 1584 28980
rect 126 28940 162 28946
rect 156 28937 162 28940
rect 810 28940 1584 28946
rect 810 28937 816 28940
rect 894 28900 900 28903
rect 126 28894 900 28900
rect 1548 28900 1554 28903
rect 1548 28894 1584 28900
rect 126 28860 138 28894
rect 1572 28860 1584 28894
rect 126 28854 900 28860
rect 894 28851 900 28854
rect 1548 28854 1584 28860
rect 1548 28851 1554 28854
rect 156 28814 162 28817
rect 126 28808 162 28814
rect 810 28814 816 28817
rect 810 28808 1584 28814
rect 126 28774 138 28808
rect 1572 28774 1584 28808
rect 126 28768 162 28774
rect 156 28765 162 28768
rect 810 28768 1584 28774
rect 810 28765 816 28768
rect 894 28728 900 28731
rect 126 28722 900 28728
rect 1548 28728 1554 28731
rect 1548 28722 1584 28728
rect 126 28688 138 28722
rect 1572 28688 1584 28722
rect 126 28682 900 28688
rect 894 28679 900 28682
rect 1548 28682 1584 28688
rect 1548 28679 1554 28682
rect 156 28642 162 28645
rect 126 28636 162 28642
rect 810 28642 816 28645
rect 810 28636 1584 28642
rect 126 28602 138 28636
rect 1572 28602 1584 28636
rect 126 28596 162 28602
rect 156 28593 162 28596
rect 810 28596 1584 28602
rect 810 28593 816 28596
rect 894 28556 900 28559
rect 126 28550 900 28556
rect 1548 28556 1554 28559
rect 1548 28550 1584 28556
rect 126 28516 138 28550
rect 1572 28516 1584 28550
rect 126 28510 900 28516
rect 894 28507 900 28510
rect 1548 28510 1584 28516
rect 1548 28507 1554 28510
rect 156 28470 162 28473
rect 126 28464 162 28470
rect 810 28470 816 28473
rect 810 28464 1584 28470
rect 126 28430 138 28464
rect 1572 28430 1584 28464
rect 126 28424 162 28430
rect 156 28421 162 28424
rect 810 28424 1584 28430
rect 810 28421 816 28424
rect 894 28384 900 28387
rect 126 28378 900 28384
rect 1548 28384 1554 28387
rect 1548 28378 1584 28384
rect 126 28344 138 28378
rect 1572 28344 1584 28378
rect 126 28338 900 28344
rect 894 28335 900 28338
rect 1548 28338 1584 28344
rect 1548 28335 1554 28338
rect 156 28298 162 28301
rect 126 28292 162 28298
rect 810 28298 816 28301
rect 810 28292 1584 28298
rect 126 28258 138 28292
rect 1572 28258 1584 28292
rect 126 28252 162 28258
rect 156 28249 162 28252
rect 810 28252 1584 28258
rect 810 28249 816 28252
rect 894 28212 900 28215
rect 126 28206 900 28212
rect 1548 28212 1554 28215
rect 1548 28206 1584 28212
rect 126 28172 138 28206
rect 1572 28172 1584 28206
rect 126 28166 900 28172
rect 894 28163 900 28166
rect 1548 28166 1584 28172
rect 1548 28163 1554 28166
rect 156 28126 162 28129
rect 126 28120 162 28126
rect 810 28126 816 28129
rect 810 28120 1584 28126
rect 126 28086 138 28120
rect 1572 28086 1584 28120
rect 126 28080 162 28086
rect 156 28077 162 28080
rect 810 28080 1584 28086
rect 810 28077 816 28080
rect 894 28040 900 28043
rect 126 28034 900 28040
rect 1548 28040 1554 28043
rect 1548 28034 1584 28040
rect 126 28000 138 28034
rect 1572 28000 1584 28034
rect 126 27994 900 28000
rect 894 27991 900 27994
rect 1548 27994 1584 28000
rect 1548 27991 1554 27994
rect 156 27954 162 27957
rect 126 27948 162 27954
rect 810 27954 816 27957
rect 810 27948 1584 27954
rect 126 27914 138 27948
rect 1572 27914 1584 27948
rect 126 27908 162 27914
rect 156 27905 162 27908
rect 810 27908 1584 27914
rect 810 27905 816 27908
rect 894 27868 900 27871
rect 126 27862 900 27868
rect 1548 27868 1554 27871
rect 1548 27862 1584 27868
rect 126 27828 138 27862
rect 1572 27828 1584 27862
rect 126 27822 900 27828
rect 894 27819 900 27822
rect 1548 27822 1584 27828
rect 1548 27819 1554 27822
rect 156 27782 162 27785
rect 126 27776 162 27782
rect 810 27782 816 27785
rect 810 27776 1584 27782
rect 126 27742 138 27776
rect 1572 27742 1584 27776
rect 126 27736 162 27742
rect 156 27733 162 27736
rect 810 27736 1584 27742
rect 810 27733 816 27736
rect 894 27696 900 27699
rect 126 27690 900 27696
rect 1548 27696 1554 27699
rect 1548 27690 1584 27696
rect 126 27656 138 27690
rect 1572 27656 1584 27690
rect 126 27650 900 27656
rect 894 27647 900 27650
rect 1548 27650 1584 27656
rect 1548 27647 1554 27650
rect 156 27610 162 27613
rect 126 27604 162 27610
rect 810 27610 816 27613
rect 810 27604 1584 27610
rect 126 27570 138 27604
rect 1572 27570 1584 27604
rect 126 27564 162 27570
rect 156 27561 162 27564
rect 810 27564 1584 27570
rect 810 27561 816 27564
rect 894 27524 900 27527
rect 126 27518 900 27524
rect 1548 27524 1554 27527
rect 1548 27518 1584 27524
rect 126 27484 138 27518
rect 1572 27484 1584 27518
rect 126 27478 900 27484
rect 894 27475 900 27478
rect 1548 27478 1584 27484
rect 1548 27475 1554 27478
rect 156 27438 162 27441
rect 126 27432 162 27438
rect 810 27438 816 27441
rect 810 27432 1584 27438
rect 126 27398 138 27432
rect 1572 27398 1584 27432
rect 126 27392 162 27398
rect 156 27389 162 27392
rect 810 27392 1584 27398
rect 810 27389 816 27392
rect 894 27352 900 27355
rect 126 27346 900 27352
rect 1548 27352 1554 27355
rect 1548 27346 1584 27352
rect 126 27312 138 27346
rect 1572 27312 1584 27346
rect 126 27306 900 27312
rect 894 27303 900 27306
rect 1548 27306 1584 27312
rect 1548 27303 1554 27306
rect 156 27266 162 27269
rect 126 27260 162 27266
rect 810 27266 816 27269
rect 810 27260 1584 27266
rect 126 27226 138 27260
rect 1572 27226 1584 27260
rect 126 27220 162 27226
rect 156 27217 162 27220
rect 810 27220 1584 27226
rect 810 27217 816 27220
rect 894 27180 900 27183
rect 126 27174 900 27180
rect 1548 27180 1554 27183
rect 1548 27174 1584 27180
rect 126 27140 138 27174
rect 1572 27140 1584 27174
rect 126 27134 900 27140
rect 894 27131 900 27134
rect 1548 27134 1584 27140
rect 1548 27131 1554 27134
rect 156 27094 162 27097
rect 126 27088 162 27094
rect 810 27094 816 27097
rect 810 27088 1584 27094
rect 126 27054 138 27088
rect 1572 27054 1584 27088
rect 126 27048 162 27054
rect 156 27045 162 27048
rect 810 27048 1584 27054
rect 810 27045 816 27048
rect 894 27008 900 27011
rect 126 27002 900 27008
rect 1548 27008 1554 27011
rect 1548 27002 1584 27008
rect 126 26968 138 27002
rect 1572 26968 1584 27002
rect 126 26962 900 26968
rect 894 26959 900 26962
rect 1548 26962 1584 26968
rect 1548 26959 1554 26962
rect 156 26922 162 26925
rect 126 26916 162 26922
rect 810 26922 816 26925
rect 810 26916 1584 26922
rect 126 26882 138 26916
rect 1572 26882 1584 26916
rect 126 26876 162 26882
rect 156 26873 162 26876
rect 810 26876 1584 26882
rect 810 26873 816 26876
rect 894 26836 900 26839
rect 126 26830 900 26836
rect 1548 26836 1554 26839
rect 1548 26830 1584 26836
rect 126 26796 138 26830
rect 1572 26796 1584 26830
rect 126 26790 900 26796
rect 894 26787 900 26790
rect 1548 26790 1584 26796
rect 1548 26787 1554 26790
rect 156 26750 162 26753
rect 126 26744 162 26750
rect 810 26750 816 26753
rect 810 26744 1584 26750
rect 126 26710 138 26744
rect 1572 26710 1584 26744
rect 126 26704 162 26710
rect 156 26701 162 26704
rect 810 26704 1584 26710
rect 810 26701 816 26704
rect 894 26664 900 26667
rect 126 26658 900 26664
rect 1548 26664 1554 26667
rect 1548 26658 1584 26664
rect 126 26624 138 26658
rect 1572 26624 1584 26658
rect 126 26618 900 26624
rect 894 26615 900 26618
rect 1548 26618 1584 26624
rect 1548 26615 1554 26618
rect 156 26578 162 26581
rect 126 26572 162 26578
rect 810 26578 816 26581
rect 810 26572 1584 26578
rect 126 26538 138 26572
rect 1572 26538 1584 26572
rect 126 26532 162 26538
rect 156 26529 162 26532
rect 810 26532 1584 26538
rect 810 26529 816 26532
rect 894 26492 900 26495
rect 126 26486 900 26492
rect 1548 26492 1554 26495
rect 1548 26486 1584 26492
rect 126 26452 138 26486
rect 1572 26452 1584 26486
rect 126 26446 900 26452
rect 894 26443 900 26446
rect 1548 26446 1584 26452
rect 1548 26443 1554 26446
rect 156 26406 162 26409
rect 126 26400 162 26406
rect 810 26406 816 26409
rect 810 26400 1584 26406
rect 126 26366 138 26400
rect 1572 26366 1584 26400
rect 126 26360 162 26366
rect 156 26357 162 26360
rect 810 26360 1584 26366
rect 810 26357 816 26360
rect 894 26320 900 26323
rect 126 26314 900 26320
rect 1548 26320 1554 26323
rect 1548 26314 1584 26320
rect 126 26280 138 26314
rect 1572 26280 1584 26314
rect 126 26274 900 26280
rect 894 26271 900 26274
rect 1548 26274 1584 26280
rect 1548 26271 1554 26274
rect 156 26234 162 26237
rect 126 26228 162 26234
rect 810 26234 816 26237
rect 810 26228 1584 26234
rect 126 26194 138 26228
rect 1572 26194 1584 26228
rect 126 26188 162 26194
rect 156 26185 162 26188
rect 810 26188 1584 26194
rect 810 26185 816 26188
rect 894 26148 900 26151
rect 126 26142 900 26148
rect 1548 26148 1554 26151
rect 1548 26142 1584 26148
rect 126 26108 138 26142
rect 1572 26108 1584 26142
rect 126 26102 900 26108
rect 894 26099 900 26102
rect 1548 26102 1584 26108
rect 1548 26099 1554 26102
rect 156 26062 162 26065
rect 126 26056 162 26062
rect 810 26062 816 26065
rect 810 26056 1584 26062
rect 126 26022 138 26056
rect 1572 26022 1584 26056
rect 126 26016 162 26022
rect 156 26013 162 26016
rect 810 26016 1584 26022
rect 810 26013 816 26016
rect 894 25976 900 25979
rect 126 25970 900 25976
rect 1548 25976 1554 25979
rect 1548 25970 1584 25976
rect 126 25936 138 25970
rect 1572 25936 1584 25970
rect 126 25930 900 25936
rect 894 25927 900 25930
rect 1548 25930 1584 25936
rect 1548 25927 1554 25930
rect 156 25890 162 25893
rect 126 25884 162 25890
rect 810 25890 816 25893
rect 810 25884 1584 25890
rect 126 25850 138 25884
rect 1572 25850 1584 25884
rect 126 25844 162 25850
rect 156 25841 162 25844
rect 810 25844 1584 25850
rect 810 25841 816 25844
rect 894 25804 900 25807
rect 126 25798 900 25804
rect 1548 25804 1554 25807
rect 1548 25798 1584 25804
rect 126 25764 138 25798
rect 1572 25764 1584 25798
rect 126 25758 900 25764
rect 894 25755 900 25758
rect 1548 25758 1584 25764
rect 1548 25755 1554 25758
rect 156 25718 162 25721
rect 126 25712 162 25718
rect 810 25718 816 25721
rect 810 25712 1584 25718
rect 126 25678 138 25712
rect 1572 25678 1584 25712
rect 126 25672 162 25678
rect 156 25669 162 25672
rect 810 25672 1584 25678
rect 810 25669 816 25672
rect 894 25632 900 25635
rect 126 25626 900 25632
rect 1548 25632 1554 25635
rect 1548 25626 1584 25632
rect 126 25592 138 25626
rect 1572 25592 1584 25626
rect 126 25586 900 25592
rect 894 25583 900 25586
rect 1548 25586 1584 25592
rect 1548 25583 1554 25586
rect 156 25546 162 25549
rect 126 25540 162 25546
rect 810 25546 816 25549
rect 810 25540 1584 25546
rect 126 25506 138 25540
rect 1572 25506 1584 25540
rect 126 25500 162 25506
rect 156 25497 162 25500
rect 810 25500 1584 25506
rect 810 25497 816 25500
rect 894 25460 900 25463
rect 126 25454 900 25460
rect 1548 25460 1554 25463
rect 1548 25454 1584 25460
rect 126 25420 138 25454
rect 1572 25420 1584 25454
rect 126 25414 900 25420
rect 894 25411 900 25414
rect 1548 25414 1584 25420
rect 1548 25411 1554 25414
rect 156 25374 162 25377
rect 126 25368 162 25374
rect 810 25374 816 25377
rect 810 25368 1584 25374
rect 126 25334 138 25368
rect 1572 25334 1584 25368
rect 126 25328 162 25334
rect 156 25325 162 25328
rect 810 25328 1584 25334
rect 810 25325 816 25328
rect 894 25288 900 25291
rect 126 25282 900 25288
rect 1548 25288 1554 25291
rect 1548 25282 1584 25288
rect 126 25248 138 25282
rect 1572 25248 1584 25282
rect 126 25242 900 25248
rect 894 25239 900 25242
rect 1548 25242 1584 25248
rect 1548 25239 1554 25242
rect 156 25202 162 25205
rect 126 25196 162 25202
rect 810 25202 816 25205
rect 810 25196 1584 25202
rect 126 25162 138 25196
rect 1572 25162 1584 25196
rect 126 25156 162 25162
rect 156 25153 162 25156
rect 810 25156 1584 25162
rect 810 25153 816 25156
rect 894 25116 900 25119
rect 126 25110 900 25116
rect 1548 25116 1554 25119
rect 1548 25110 1584 25116
rect 126 25076 138 25110
rect 1572 25076 1584 25110
rect 126 25070 900 25076
rect 894 25067 900 25070
rect 1548 25070 1584 25076
rect 1548 25067 1554 25070
rect 156 25030 162 25033
rect 126 25024 162 25030
rect 810 25030 816 25033
rect 810 25024 1584 25030
rect 126 24990 138 25024
rect 1572 24990 1584 25024
rect 126 24984 162 24990
rect 156 24981 162 24984
rect 810 24984 1584 24990
rect 810 24981 816 24984
rect 894 24944 900 24947
rect 126 24938 900 24944
rect 1548 24944 1554 24947
rect 1548 24938 1584 24944
rect 126 24904 138 24938
rect 1572 24904 1584 24938
rect 126 24898 900 24904
rect 894 24895 900 24898
rect 1548 24898 1584 24904
rect 1548 24895 1554 24898
rect 156 24858 162 24861
rect 126 24852 162 24858
rect 810 24858 816 24861
rect 810 24852 1584 24858
rect 126 24818 138 24852
rect 1572 24818 1584 24852
rect 126 24812 162 24818
rect 156 24809 162 24812
rect 810 24812 1584 24818
rect 810 24809 816 24812
rect 894 24772 900 24775
rect 126 24766 900 24772
rect 1548 24772 1554 24775
rect 1548 24766 1584 24772
rect 126 24732 138 24766
rect 1572 24732 1584 24766
rect 126 24726 900 24732
rect 894 24723 900 24726
rect 1548 24726 1584 24732
rect 1548 24723 1554 24726
rect 156 24686 162 24689
rect 126 24680 162 24686
rect 810 24686 816 24689
rect 810 24680 1584 24686
rect 126 24646 138 24680
rect 1572 24646 1584 24680
rect 126 24640 162 24646
rect 156 24637 162 24640
rect 810 24640 1584 24646
rect 810 24637 816 24640
rect 894 24600 900 24603
rect 126 24594 900 24600
rect 1548 24600 1554 24603
rect 1548 24594 1584 24600
rect 126 24560 138 24594
rect 1572 24560 1584 24594
rect 126 24554 900 24560
rect 894 24551 900 24554
rect 1548 24554 1584 24560
rect 1548 24551 1554 24554
rect 156 24514 162 24517
rect 126 24508 162 24514
rect 810 24514 816 24517
rect 810 24508 1584 24514
rect 126 24474 138 24508
rect 1572 24474 1584 24508
rect 126 24468 162 24474
rect 156 24465 162 24468
rect 810 24468 1584 24474
rect 810 24465 816 24468
rect 894 24428 900 24431
rect 126 24422 900 24428
rect 1548 24428 1554 24431
rect 1548 24422 1584 24428
rect 126 24388 138 24422
rect 1572 24388 1584 24422
rect 126 24382 900 24388
rect 894 24379 900 24382
rect 1548 24382 1584 24388
rect 1548 24379 1554 24382
rect 156 24342 162 24345
rect 126 24336 162 24342
rect 810 24342 816 24345
rect 810 24336 1584 24342
rect 126 24302 138 24336
rect 1572 24302 1584 24336
rect 126 24296 162 24302
rect 156 24293 162 24296
rect 810 24296 1584 24302
rect 810 24293 816 24296
rect 894 24256 900 24259
rect 126 24250 900 24256
rect 1548 24256 1554 24259
rect 1548 24250 1584 24256
rect 126 24216 138 24250
rect 1572 24216 1584 24250
rect 126 24210 900 24216
rect 894 24207 900 24210
rect 1548 24210 1584 24216
rect 1548 24207 1554 24210
rect 156 24170 162 24173
rect 126 24164 162 24170
rect 810 24170 816 24173
rect 810 24164 1584 24170
rect 126 24130 138 24164
rect 1572 24130 1584 24164
rect 126 24124 162 24130
rect 156 24121 162 24124
rect 810 24124 1584 24130
rect 810 24121 816 24124
rect 894 24084 900 24087
rect 126 24078 900 24084
rect 1548 24084 1554 24087
rect 1548 24078 1584 24084
rect 126 24044 138 24078
rect 1572 24044 1584 24078
rect 126 24038 900 24044
rect 894 24035 900 24038
rect 1548 24038 1584 24044
rect 1548 24035 1554 24038
rect 156 23998 162 24001
rect 126 23992 162 23998
rect 810 23998 816 24001
rect 810 23992 1584 23998
rect 126 23958 138 23992
rect 1572 23958 1584 23992
rect 126 23952 162 23958
rect 156 23949 162 23952
rect 810 23952 1584 23958
rect 810 23949 816 23952
rect 894 23912 900 23915
rect 126 23906 900 23912
rect 1548 23912 1554 23915
rect 1548 23906 1584 23912
rect 126 23872 138 23906
rect 1572 23872 1584 23906
rect 126 23866 900 23872
rect 894 23863 900 23866
rect 1548 23866 1584 23872
rect 1548 23863 1554 23866
rect 156 23826 162 23829
rect 126 23820 162 23826
rect 810 23826 816 23829
rect 810 23820 1584 23826
rect 126 23786 138 23820
rect 1572 23786 1584 23820
rect 126 23780 162 23786
rect 156 23777 162 23780
rect 810 23780 1584 23786
rect 810 23777 816 23780
rect 894 23740 900 23743
rect 126 23734 900 23740
rect 1548 23740 1554 23743
rect 1548 23734 1584 23740
rect 126 23700 138 23734
rect 1572 23700 1584 23734
rect 126 23694 900 23700
rect 894 23691 900 23694
rect 1548 23694 1584 23700
rect 1548 23691 1554 23694
rect 156 23654 162 23657
rect 126 23648 162 23654
rect 810 23654 816 23657
rect 810 23648 1584 23654
rect 126 23614 138 23648
rect 1572 23614 1584 23648
rect 126 23608 162 23614
rect 156 23605 162 23608
rect 810 23608 1584 23614
rect 810 23605 816 23608
rect 894 23568 900 23571
rect 126 23562 900 23568
rect 1548 23568 1554 23571
rect 1548 23562 1584 23568
rect 126 23528 138 23562
rect 1572 23528 1584 23562
rect 126 23522 900 23528
rect 894 23519 900 23522
rect 1548 23522 1584 23528
rect 1548 23519 1554 23522
rect 156 23482 162 23485
rect 126 23476 162 23482
rect 810 23482 816 23485
rect 810 23476 1584 23482
rect 126 23442 138 23476
rect 1572 23442 1584 23476
rect 126 23436 162 23442
rect 156 23433 162 23436
rect 810 23436 1584 23442
rect 810 23433 816 23436
rect 894 23396 900 23399
rect 126 23390 900 23396
rect 1548 23396 1554 23399
rect 1548 23390 1584 23396
rect 126 23356 138 23390
rect 1572 23356 1584 23390
rect 126 23350 900 23356
rect 894 23347 900 23350
rect 1548 23350 1584 23356
rect 1548 23347 1554 23350
rect 156 23310 162 23313
rect 126 23304 162 23310
rect 810 23310 816 23313
rect 810 23304 1584 23310
rect 126 23270 138 23304
rect 1572 23270 1584 23304
rect 126 23264 162 23270
rect 156 23261 162 23264
rect 810 23264 1584 23270
rect 810 23261 816 23264
rect 894 23224 900 23227
rect 126 23218 900 23224
rect 1548 23224 1554 23227
rect 1548 23218 1584 23224
rect 126 23184 138 23218
rect 1572 23184 1584 23218
rect 126 23178 900 23184
rect 894 23175 900 23178
rect 1548 23178 1584 23184
rect 1548 23175 1554 23178
rect 156 23138 162 23141
rect 126 23132 162 23138
rect 810 23138 816 23141
rect 810 23132 1584 23138
rect 126 23098 138 23132
rect 1572 23098 1584 23132
rect 126 23092 162 23098
rect 156 23089 162 23092
rect 810 23092 1584 23098
rect 810 23089 816 23092
rect 894 23052 900 23055
rect 126 23046 900 23052
rect 1548 23052 1554 23055
rect 1548 23046 1584 23052
rect 126 23012 138 23046
rect 1572 23012 1584 23046
rect 126 23006 900 23012
rect 894 23003 900 23006
rect 1548 23006 1584 23012
rect 1548 23003 1554 23006
rect 156 22966 162 22969
rect 126 22960 162 22966
rect 810 22966 816 22969
rect 810 22960 1584 22966
rect 126 22926 138 22960
rect 1572 22926 1584 22960
rect 126 22920 162 22926
rect 156 22917 162 22920
rect 810 22920 1584 22926
rect 810 22917 816 22920
rect 894 22880 900 22883
rect 126 22874 900 22880
rect 1548 22880 1554 22883
rect 1548 22874 1584 22880
rect 126 22840 138 22874
rect 1572 22840 1584 22874
rect 126 22834 900 22840
rect 894 22831 900 22834
rect 1548 22834 1584 22840
rect 1548 22831 1554 22834
rect 156 22794 162 22797
rect 126 22788 162 22794
rect 810 22794 816 22797
rect 810 22788 1584 22794
rect 126 22754 138 22788
rect 1572 22754 1584 22788
rect 126 22748 162 22754
rect 156 22745 162 22748
rect 810 22748 1584 22754
rect 810 22745 816 22748
rect 894 22708 900 22711
rect 126 22702 900 22708
rect 1548 22708 1554 22711
rect 1548 22702 1584 22708
rect 126 22668 138 22702
rect 1572 22668 1584 22702
rect 126 22662 900 22668
rect 894 22659 900 22662
rect 1548 22662 1584 22668
rect 1548 22659 1554 22662
rect 156 22622 162 22625
rect 126 22616 162 22622
rect 810 22622 816 22625
rect 810 22616 1584 22622
rect 126 22582 138 22616
rect 1572 22582 1584 22616
rect 126 22576 162 22582
rect 156 22573 162 22576
rect 810 22576 1584 22582
rect 810 22573 816 22576
rect 894 22536 900 22539
rect 126 22530 900 22536
rect 1548 22536 1554 22539
rect 1548 22530 1584 22536
rect 126 22496 138 22530
rect 1572 22496 1584 22530
rect 126 22490 900 22496
rect 894 22487 900 22490
rect 1548 22490 1584 22496
rect 1548 22487 1554 22490
rect 156 22450 162 22453
rect 126 22444 162 22450
rect 810 22450 816 22453
rect 810 22444 1584 22450
rect 126 22410 138 22444
rect 1572 22410 1584 22444
rect 126 22404 162 22410
rect 156 22401 162 22404
rect 810 22404 1584 22410
rect 810 22401 816 22404
rect 894 22364 900 22367
rect 126 22358 900 22364
rect 1548 22364 1554 22367
rect 1548 22358 1584 22364
rect 126 22324 138 22358
rect 1572 22324 1584 22358
rect 126 22318 900 22324
rect 894 22315 900 22318
rect 1548 22318 1584 22324
rect 1548 22315 1554 22318
rect 156 22278 162 22281
rect 126 22272 162 22278
rect 810 22278 816 22281
rect 810 22272 1584 22278
rect 126 22238 138 22272
rect 1572 22238 1584 22272
rect 126 22232 162 22238
rect 156 22229 162 22232
rect 810 22232 1584 22238
rect 810 22229 816 22232
rect 894 22192 900 22195
rect 126 22186 900 22192
rect 1548 22192 1554 22195
rect 1548 22186 1584 22192
rect 126 22152 138 22186
rect 1572 22152 1584 22186
rect 126 22146 900 22152
rect 894 22143 900 22146
rect 1548 22146 1584 22152
rect 1548 22143 1554 22146
rect 156 22106 162 22109
rect 126 22100 162 22106
rect 810 22106 816 22109
rect 810 22100 1584 22106
rect 126 22066 138 22100
rect 1572 22066 1584 22100
rect 126 22060 162 22066
rect 156 22057 162 22060
rect 810 22060 1584 22066
rect 810 22057 816 22060
rect 894 22020 900 22023
rect 126 22014 900 22020
rect 1548 22020 1554 22023
rect 1548 22014 1584 22020
rect 126 21980 138 22014
rect 1572 21980 1584 22014
rect 126 21974 900 21980
rect 894 21971 900 21974
rect 1548 21974 1584 21980
rect 1548 21971 1554 21974
rect 156 21934 162 21937
rect 126 21928 162 21934
rect 810 21934 816 21937
rect 810 21928 1584 21934
rect 126 21894 138 21928
rect 1572 21894 1584 21928
rect 126 21888 162 21894
rect 156 21885 162 21888
rect 810 21888 1584 21894
rect 810 21885 816 21888
rect 894 21848 900 21851
rect 126 21842 900 21848
rect 1548 21848 1554 21851
rect 1548 21842 1584 21848
rect 126 21808 138 21842
rect 1572 21808 1584 21842
rect 126 21802 900 21808
rect 894 21799 900 21802
rect 1548 21802 1584 21808
rect 1548 21799 1554 21802
rect 156 21762 162 21765
rect 126 21756 162 21762
rect 810 21762 816 21765
rect 810 21756 1584 21762
rect 126 21722 138 21756
rect 1572 21722 1584 21756
rect 126 21716 162 21722
rect 156 21713 162 21716
rect 810 21716 1584 21722
rect 810 21713 816 21716
rect 894 21676 900 21679
rect 126 21670 900 21676
rect 1548 21676 1554 21679
rect 1548 21670 1584 21676
rect 126 21636 138 21670
rect 1572 21636 1584 21670
rect 126 21630 900 21636
rect 894 21627 900 21630
rect 1548 21630 1584 21636
rect 1548 21627 1554 21630
rect 156 21590 162 21593
rect 126 21584 162 21590
rect 810 21590 816 21593
rect 810 21584 1584 21590
rect 126 21550 138 21584
rect 1572 21550 1584 21584
rect 126 21544 162 21550
rect 156 21541 162 21544
rect 810 21544 1584 21550
rect 810 21541 816 21544
rect 894 21504 900 21507
rect 126 21498 900 21504
rect 1548 21504 1554 21507
rect 1548 21498 1584 21504
rect 126 21464 138 21498
rect 1572 21464 1584 21498
rect 126 21458 900 21464
rect 894 21455 900 21458
rect 1548 21458 1584 21464
rect 1548 21455 1554 21458
rect 156 21418 162 21421
rect 126 21412 162 21418
rect 810 21418 816 21421
rect 810 21412 1584 21418
rect 126 21378 138 21412
rect 1572 21378 1584 21412
rect 126 21372 162 21378
rect 156 21369 162 21372
rect 810 21372 1584 21378
rect 810 21369 816 21372
rect 894 21332 900 21335
rect 126 21326 900 21332
rect 1548 21332 1554 21335
rect 1548 21326 1584 21332
rect 126 21292 138 21326
rect 1572 21292 1584 21326
rect 126 21286 900 21292
rect 894 21283 900 21286
rect 1548 21286 1584 21292
rect 1548 21283 1554 21286
rect 156 21246 162 21249
rect 126 21240 162 21246
rect 810 21246 816 21249
rect 810 21240 1584 21246
rect 126 21206 138 21240
rect 1572 21206 1584 21240
rect 126 21200 162 21206
rect 156 21197 162 21200
rect 810 21200 1584 21206
rect 810 21197 816 21200
rect 894 21160 900 21163
rect 126 21154 900 21160
rect 1548 21160 1554 21163
rect 1548 21154 1584 21160
rect 126 21120 138 21154
rect 1572 21120 1584 21154
rect 126 21114 900 21120
rect 894 21111 900 21114
rect 1548 21114 1584 21120
rect 1548 21111 1554 21114
rect 156 21074 162 21077
rect 126 21068 162 21074
rect 810 21074 816 21077
rect 810 21068 1584 21074
rect 126 21034 138 21068
rect 1572 21034 1584 21068
rect 126 21028 162 21034
rect 156 21025 162 21028
rect 810 21028 1584 21034
rect 810 21025 816 21028
rect 894 20988 900 20991
rect 126 20982 900 20988
rect 1548 20988 1554 20991
rect 1548 20982 1584 20988
rect 126 20948 138 20982
rect 1572 20948 1584 20982
rect 126 20942 900 20948
rect 894 20939 900 20942
rect 1548 20942 1584 20948
rect 1548 20939 1554 20942
rect 156 20902 162 20905
rect 126 20896 162 20902
rect 810 20902 816 20905
rect 810 20896 1584 20902
rect 126 20862 138 20896
rect 1572 20862 1584 20896
rect 126 20856 162 20862
rect 156 20853 162 20856
rect 810 20856 1584 20862
rect 810 20853 816 20856
rect 894 20816 900 20819
rect 126 20810 900 20816
rect 1548 20816 1554 20819
rect 1548 20810 1584 20816
rect 126 20776 138 20810
rect 1572 20776 1584 20810
rect 126 20770 900 20776
rect 894 20767 900 20770
rect 1548 20770 1584 20776
rect 1548 20767 1554 20770
rect 156 20730 162 20733
rect 126 20724 162 20730
rect 810 20730 816 20733
rect 810 20724 1584 20730
rect 126 20690 138 20724
rect 1572 20690 1584 20724
rect 126 20684 162 20690
rect 156 20681 162 20684
rect 810 20684 1584 20690
rect 810 20681 816 20684
rect 894 20644 900 20647
rect 126 20638 900 20644
rect 1548 20644 1554 20647
rect 1548 20638 1584 20644
rect 126 20604 138 20638
rect 1572 20604 1584 20638
rect 126 20598 900 20604
rect 894 20595 900 20598
rect 1548 20598 1584 20604
rect 1548 20595 1554 20598
rect 156 20558 162 20561
rect 126 20552 162 20558
rect 810 20558 816 20561
rect 810 20552 1584 20558
rect 126 20518 138 20552
rect 1572 20518 1584 20552
rect 126 20512 162 20518
rect 156 20509 162 20512
rect 810 20512 1584 20518
rect 810 20509 816 20512
rect 894 20472 900 20475
rect 126 20466 900 20472
rect 1548 20472 1554 20475
rect 1548 20466 1584 20472
rect 126 20432 138 20466
rect 1572 20432 1584 20466
rect 126 20426 900 20432
rect 894 20423 900 20426
rect 1548 20426 1584 20432
rect 1548 20423 1554 20426
rect 156 20386 162 20389
rect 126 20380 162 20386
rect 810 20386 816 20389
rect 810 20380 1584 20386
rect 126 20346 138 20380
rect 1572 20346 1584 20380
rect 126 20340 162 20346
rect 156 20337 162 20340
rect 810 20340 1584 20346
rect 810 20337 816 20340
rect 894 20300 900 20303
rect 126 20294 900 20300
rect 1548 20300 1554 20303
rect 1548 20294 1584 20300
rect 126 20260 138 20294
rect 1572 20260 1584 20294
rect 126 20254 900 20260
rect 894 20251 900 20254
rect 1548 20254 1584 20260
rect 1548 20251 1554 20254
rect 156 20214 162 20217
rect 126 20208 162 20214
rect 810 20214 816 20217
rect 810 20208 1584 20214
rect 126 20174 138 20208
rect 1572 20174 1584 20208
rect 126 20168 162 20174
rect 156 20165 162 20168
rect 810 20168 1584 20174
rect 810 20165 816 20168
rect 894 20128 900 20131
rect 126 20122 900 20128
rect 1548 20128 1554 20131
rect 1548 20122 1584 20128
rect 126 20088 138 20122
rect 1572 20088 1584 20122
rect 126 20082 900 20088
rect 894 20079 900 20082
rect 1548 20082 1584 20088
rect 1548 20079 1554 20082
rect 156 20042 162 20045
rect 126 20036 162 20042
rect 810 20042 816 20045
rect 810 20036 1584 20042
rect 126 20002 138 20036
rect 1572 20002 1584 20036
rect 126 19996 162 20002
rect 156 19993 162 19996
rect 810 19996 1584 20002
rect 810 19993 816 19996
rect 894 19956 900 19959
rect 126 19950 900 19956
rect 1548 19956 1554 19959
rect 1548 19950 1584 19956
rect 126 19916 138 19950
rect 1572 19916 1584 19950
rect 126 19910 900 19916
rect 894 19907 900 19910
rect 1548 19910 1584 19916
rect 1548 19907 1554 19910
rect 156 19870 162 19873
rect 126 19864 162 19870
rect 810 19870 816 19873
rect 810 19864 1584 19870
rect 126 19830 138 19864
rect 1572 19830 1584 19864
rect 126 19824 162 19830
rect 156 19821 162 19824
rect 810 19824 1584 19830
rect 810 19821 816 19824
rect 894 19784 900 19787
rect 126 19778 900 19784
rect 1548 19784 1554 19787
rect 1548 19778 1584 19784
rect 126 19744 138 19778
rect 1572 19744 1584 19778
rect 126 19738 900 19744
rect 894 19735 900 19738
rect 1548 19738 1584 19744
rect 1548 19735 1554 19738
rect 156 19698 162 19701
rect 126 19692 162 19698
rect 810 19698 816 19701
rect 810 19692 1584 19698
rect 126 19658 138 19692
rect 1572 19658 1584 19692
rect 126 19652 162 19658
rect 156 19649 162 19652
rect 810 19652 1584 19658
rect 810 19649 816 19652
rect 894 19612 900 19615
rect 126 19606 900 19612
rect 1548 19612 1554 19615
rect 1548 19606 1584 19612
rect 126 19572 138 19606
rect 1572 19572 1584 19606
rect 126 19566 900 19572
rect 894 19563 900 19566
rect 1548 19566 1584 19572
rect 1548 19563 1554 19566
rect 156 19526 162 19529
rect 126 19520 162 19526
rect 810 19526 816 19529
rect 810 19520 1584 19526
rect 126 19486 138 19520
rect 1572 19486 1584 19520
rect 126 19480 162 19486
rect 156 19477 162 19480
rect 810 19480 1584 19486
rect 810 19477 816 19480
rect 894 19440 900 19443
rect 126 19434 900 19440
rect 1548 19440 1554 19443
rect 1548 19434 1584 19440
rect 126 19400 138 19434
rect 1572 19400 1584 19434
rect 126 19394 900 19400
rect 894 19391 900 19394
rect 1548 19394 1584 19400
rect 1548 19391 1554 19394
rect 156 19354 162 19357
rect 126 19348 162 19354
rect 810 19354 816 19357
rect 810 19348 1584 19354
rect 126 19314 138 19348
rect 1572 19314 1584 19348
rect 126 19308 162 19314
rect 156 19305 162 19308
rect 810 19308 1584 19314
rect 810 19305 816 19308
rect 894 19268 900 19271
rect 126 19262 900 19268
rect 1548 19268 1554 19271
rect 1548 19262 1584 19268
rect 126 19228 138 19262
rect 1572 19228 1584 19262
rect 126 19222 900 19228
rect 894 19219 900 19222
rect 1548 19222 1584 19228
rect 1548 19219 1554 19222
rect 156 19182 162 19185
rect 126 19176 162 19182
rect 810 19182 816 19185
rect 810 19176 1584 19182
rect 126 19142 138 19176
rect 1572 19142 1584 19176
rect 126 19136 162 19142
rect 156 19133 162 19136
rect 810 19136 1584 19142
rect 810 19133 816 19136
rect 894 19096 900 19099
rect 126 19090 900 19096
rect 1548 19096 1554 19099
rect 1548 19090 1584 19096
rect 126 19056 138 19090
rect 1572 19056 1584 19090
rect 126 19050 900 19056
rect 894 19047 900 19050
rect 1548 19050 1584 19056
rect 1548 19047 1554 19050
rect 156 19010 162 19013
rect 126 19004 162 19010
rect 810 19010 816 19013
rect 810 19004 1584 19010
rect 126 18970 138 19004
rect 1572 18970 1584 19004
rect 126 18964 162 18970
rect 156 18961 162 18964
rect 810 18964 1584 18970
rect 810 18961 816 18964
rect 894 18924 900 18927
rect 126 18918 900 18924
rect 1548 18924 1554 18927
rect 1548 18918 1584 18924
rect 126 18884 138 18918
rect 1572 18884 1584 18918
rect 126 18878 900 18884
rect 894 18875 900 18878
rect 1548 18878 1584 18884
rect 1548 18875 1554 18878
rect 156 18838 162 18841
rect 126 18832 162 18838
rect 810 18838 816 18841
rect 810 18832 1584 18838
rect 126 18798 138 18832
rect 1572 18798 1584 18832
rect 126 18792 162 18798
rect 156 18789 162 18792
rect 810 18792 1584 18798
rect 810 18789 816 18792
rect 894 18752 900 18755
rect 126 18746 900 18752
rect 1548 18752 1554 18755
rect 1548 18746 1584 18752
rect 126 18712 138 18746
rect 1572 18712 1584 18746
rect 126 18706 900 18712
rect 894 18703 900 18706
rect 1548 18706 1584 18712
rect 1548 18703 1554 18706
rect 156 18666 162 18669
rect 126 18660 162 18666
rect 810 18666 816 18669
rect 810 18660 1584 18666
rect 126 18626 138 18660
rect 1572 18626 1584 18660
rect 126 18620 162 18626
rect 156 18617 162 18620
rect 810 18620 1584 18626
rect 810 18617 816 18620
rect 894 18580 900 18583
rect 126 18574 900 18580
rect 1548 18580 1554 18583
rect 1548 18574 1584 18580
rect 126 18540 138 18574
rect 1572 18540 1584 18574
rect 126 18534 900 18540
rect 894 18531 900 18534
rect 1548 18534 1584 18540
rect 1548 18531 1554 18534
rect 156 18494 162 18497
rect 126 18488 162 18494
rect 810 18494 816 18497
rect 810 18488 1584 18494
rect 126 18454 138 18488
rect 1572 18454 1584 18488
rect 126 18448 162 18454
rect 156 18445 162 18448
rect 810 18448 1584 18454
rect 810 18445 816 18448
rect 894 18408 900 18411
rect 126 18402 900 18408
rect 1548 18408 1554 18411
rect 1548 18402 1584 18408
rect 126 18368 138 18402
rect 1572 18368 1584 18402
rect 126 18362 900 18368
rect 894 18359 900 18362
rect 1548 18362 1584 18368
rect 1548 18359 1554 18362
rect 156 18322 162 18325
rect 126 18316 162 18322
rect 810 18322 816 18325
rect 810 18316 1584 18322
rect 126 18282 138 18316
rect 1572 18282 1584 18316
rect 126 18276 162 18282
rect 156 18273 162 18276
rect 810 18276 1584 18282
rect 810 18273 816 18276
rect 894 18236 900 18239
rect 126 18230 900 18236
rect 1548 18236 1554 18239
rect 1548 18230 1584 18236
rect 126 18196 138 18230
rect 1572 18196 1584 18230
rect 126 18190 900 18196
rect 894 18187 900 18190
rect 1548 18190 1584 18196
rect 1548 18187 1554 18190
rect 156 18150 162 18153
rect 126 18144 162 18150
rect 810 18150 816 18153
rect 810 18144 1584 18150
rect 126 18110 138 18144
rect 1572 18110 1584 18144
rect 126 18104 162 18110
rect 156 18101 162 18104
rect 810 18104 1584 18110
rect 810 18101 816 18104
rect 894 18064 900 18067
rect 126 18058 900 18064
rect 1548 18064 1554 18067
rect 1548 18058 1584 18064
rect 126 18024 138 18058
rect 1572 18024 1584 18058
rect 126 18018 900 18024
rect 894 18015 900 18018
rect 1548 18018 1584 18024
rect 1548 18015 1554 18018
rect 156 17978 162 17981
rect 126 17972 162 17978
rect 810 17978 816 17981
rect 810 17972 1584 17978
rect 126 17938 138 17972
rect 1572 17938 1584 17972
rect 126 17932 162 17938
rect 156 17929 162 17932
rect 810 17932 1584 17938
rect 810 17929 816 17932
rect 894 17892 900 17895
rect 126 17886 900 17892
rect 1548 17892 1554 17895
rect 1548 17886 1584 17892
rect 126 17852 138 17886
rect 1572 17852 1584 17886
rect 126 17846 900 17852
rect 894 17843 900 17846
rect 1548 17846 1584 17852
rect 1548 17843 1554 17846
rect 156 17806 162 17809
rect 126 17800 162 17806
rect 810 17806 816 17809
rect 810 17800 1584 17806
rect 126 17766 138 17800
rect 1572 17766 1584 17800
rect 126 17760 162 17766
rect 156 17757 162 17760
rect 810 17760 1584 17766
rect 810 17757 816 17760
rect 894 17720 900 17723
rect 126 17714 900 17720
rect 1548 17720 1554 17723
rect 1548 17714 1584 17720
rect 126 17680 138 17714
rect 1572 17680 1584 17714
rect 126 17674 900 17680
rect 894 17671 900 17674
rect 1548 17674 1584 17680
rect 1548 17671 1554 17674
rect 156 17634 162 17637
rect 126 17628 162 17634
rect 810 17634 816 17637
rect 810 17628 1584 17634
rect 126 17594 138 17628
rect 1572 17594 1584 17628
rect 126 17588 162 17594
rect 156 17585 162 17588
rect 810 17588 1584 17594
rect 810 17585 816 17588
rect 894 17548 900 17551
rect 126 17542 900 17548
rect 1548 17548 1554 17551
rect 1548 17542 1584 17548
rect 126 17508 138 17542
rect 1572 17508 1584 17542
rect 126 17502 900 17508
rect 894 17499 900 17502
rect 1548 17502 1584 17508
rect 1548 17499 1554 17502
rect 156 17462 162 17465
rect 126 17456 162 17462
rect 810 17462 816 17465
rect 810 17456 1584 17462
rect 126 17422 138 17456
rect 1572 17422 1584 17456
rect 126 17416 162 17422
rect 156 17413 162 17416
rect 810 17416 1584 17422
rect 810 17413 816 17416
rect 894 17376 900 17379
rect 126 17370 900 17376
rect 1548 17376 1554 17379
rect 1548 17370 1584 17376
rect 126 17336 138 17370
rect 1572 17336 1584 17370
rect 126 17330 900 17336
rect 894 17327 900 17330
rect 1548 17330 1584 17336
rect 1548 17327 1554 17330
rect 156 17290 162 17293
rect 126 17284 162 17290
rect 810 17290 816 17293
rect 810 17284 1584 17290
rect 126 17250 138 17284
rect 1572 17250 1584 17284
rect 126 17244 162 17250
rect 156 17241 162 17244
rect 810 17244 1584 17250
rect 810 17241 816 17244
rect 894 17204 900 17207
rect 126 17198 900 17204
rect 1548 17204 1554 17207
rect 1548 17198 1584 17204
rect 126 17164 138 17198
rect 1572 17164 1584 17198
rect 126 17158 900 17164
rect 894 17155 900 17158
rect 1548 17158 1584 17164
rect 1548 17155 1554 17158
rect 156 17118 162 17121
rect 126 17112 162 17118
rect 810 17118 816 17121
rect 810 17112 1584 17118
rect 126 17078 138 17112
rect 1572 17078 1584 17112
rect 126 17072 162 17078
rect 156 17069 162 17072
rect 810 17072 1584 17078
rect 810 17069 816 17072
rect 894 17032 900 17035
rect 126 17026 900 17032
rect 1548 17032 1554 17035
rect 1548 17026 1584 17032
rect 126 16992 138 17026
rect 1572 16992 1584 17026
rect 126 16986 900 16992
rect 894 16983 900 16986
rect 1548 16986 1584 16992
rect 1548 16983 1554 16986
rect 156 16946 162 16949
rect 126 16940 162 16946
rect 810 16946 816 16949
rect 810 16940 1584 16946
rect 126 16906 138 16940
rect 1572 16906 1584 16940
rect 126 16900 162 16906
rect 156 16897 162 16900
rect 810 16900 1584 16906
rect 810 16897 816 16900
rect 894 16860 900 16863
rect 126 16854 900 16860
rect 1548 16860 1554 16863
rect 1548 16854 1584 16860
rect 126 16820 138 16854
rect 1572 16820 1584 16854
rect 126 16814 900 16820
rect 894 16811 900 16814
rect 1548 16814 1584 16820
rect 1548 16811 1554 16814
rect 156 16774 162 16777
rect 126 16768 162 16774
rect 810 16774 816 16777
rect 810 16768 1584 16774
rect 126 16734 138 16768
rect 1572 16734 1584 16768
rect 126 16728 162 16734
rect 156 16725 162 16728
rect 810 16728 1584 16734
rect 810 16725 816 16728
rect 894 16688 900 16691
rect 126 16682 900 16688
rect 1548 16688 1554 16691
rect 1548 16682 1584 16688
rect 126 16648 138 16682
rect 1572 16648 1584 16682
rect 126 16642 900 16648
rect 894 16639 900 16642
rect 1548 16642 1584 16648
rect 1548 16639 1554 16642
rect 156 16602 162 16605
rect 126 16596 162 16602
rect 810 16602 816 16605
rect 810 16596 1584 16602
rect 126 16562 138 16596
rect 1572 16562 1584 16596
rect 126 16556 162 16562
rect 156 16553 162 16556
rect 810 16556 1584 16562
rect 810 16553 816 16556
rect 894 16516 900 16519
rect 126 16510 900 16516
rect 1548 16516 1554 16519
rect 1548 16510 1584 16516
rect 126 16476 138 16510
rect 1572 16476 1584 16510
rect 126 16470 900 16476
rect 894 16467 900 16470
rect 1548 16470 1584 16476
rect 1548 16467 1554 16470
rect 156 16430 162 16433
rect 126 16424 162 16430
rect 810 16430 816 16433
rect 810 16424 1584 16430
rect 126 16390 138 16424
rect 1572 16390 1584 16424
rect 126 16384 162 16390
rect 156 16381 162 16384
rect 810 16384 1584 16390
rect 810 16381 816 16384
rect 894 16344 900 16347
rect 126 16338 900 16344
rect 1548 16344 1554 16347
rect 1548 16338 1584 16344
rect 126 16304 138 16338
rect 1572 16304 1584 16338
rect 126 16298 900 16304
rect 894 16295 900 16298
rect 1548 16298 1584 16304
rect 1548 16295 1554 16298
rect 156 16258 162 16261
rect 126 16252 162 16258
rect 810 16258 816 16261
rect 810 16252 1584 16258
rect 126 16218 138 16252
rect 1572 16218 1584 16252
rect 126 16212 162 16218
rect 156 16209 162 16212
rect 810 16212 1584 16218
rect 810 16209 816 16212
rect 894 16172 900 16175
rect 126 16166 900 16172
rect 1548 16172 1554 16175
rect 1548 16166 1584 16172
rect 126 16132 138 16166
rect 1572 16132 1584 16166
rect 126 16126 900 16132
rect 894 16123 900 16126
rect 1548 16126 1584 16132
rect 1548 16123 1554 16126
rect 156 16086 162 16089
rect 126 16080 162 16086
rect 810 16086 816 16089
rect 810 16080 1584 16086
rect 126 16046 138 16080
rect 1572 16046 1584 16080
rect 126 16040 162 16046
rect 156 16037 162 16040
rect 810 16040 1584 16046
rect 810 16037 816 16040
rect 894 16000 900 16003
rect 126 15994 900 16000
rect 1548 16000 1554 16003
rect 1548 15994 1584 16000
rect 126 15960 138 15994
rect 1572 15960 1584 15994
rect 126 15954 900 15960
rect 894 15951 900 15954
rect 1548 15954 1584 15960
rect 1548 15951 1554 15954
rect 156 15914 162 15917
rect 126 15908 162 15914
rect 810 15914 816 15917
rect 810 15908 1584 15914
rect 126 15874 138 15908
rect 1572 15874 1584 15908
rect 126 15868 162 15874
rect 156 15865 162 15868
rect 810 15868 1584 15874
rect 810 15865 816 15868
rect 894 15828 900 15831
rect 126 15822 900 15828
rect 1548 15828 1554 15831
rect 1548 15822 1584 15828
rect 126 15788 138 15822
rect 1572 15788 1584 15822
rect 126 15782 900 15788
rect 894 15779 900 15782
rect 1548 15782 1584 15788
rect 1548 15779 1554 15782
rect 156 15742 162 15745
rect 126 15736 162 15742
rect 810 15742 816 15745
rect 810 15736 1584 15742
rect 126 15702 138 15736
rect 1572 15702 1584 15736
rect 126 15696 162 15702
rect 156 15693 162 15696
rect 810 15696 1584 15702
rect 810 15693 816 15696
rect 894 15656 900 15659
rect 126 15650 900 15656
rect 1548 15656 1554 15659
rect 1548 15650 1584 15656
rect 126 15616 138 15650
rect 1572 15616 1584 15650
rect 126 15610 900 15616
rect 894 15607 900 15610
rect 1548 15610 1584 15616
rect 1548 15607 1554 15610
rect 156 15570 162 15573
rect 126 15564 162 15570
rect 810 15570 816 15573
rect 810 15564 1584 15570
rect 126 15530 138 15564
rect 1572 15530 1584 15564
rect 126 15524 162 15530
rect 156 15521 162 15524
rect 810 15524 1584 15530
rect 810 15521 816 15524
rect 894 15484 900 15487
rect 126 15478 900 15484
rect 1548 15484 1554 15487
rect 1548 15478 1584 15484
rect 126 15444 138 15478
rect 1572 15444 1584 15478
rect 126 15438 900 15444
rect 894 15435 900 15438
rect 1548 15438 1584 15444
rect 1548 15435 1554 15438
rect 156 15398 162 15401
rect 126 15392 162 15398
rect 810 15398 816 15401
rect 810 15392 1584 15398
rect 126 15358 138 15392
rect 1572 15358 1584 15392
rect 126 15352 162 15358
rect 156 15349 162 15352
rect 810 15352 1584 15358
rect 810 15349 816 15352
rect 894 15312 900 15315
rect 126 15306 900 15312
rect 1548 15312 1554 15315
rect 1548 15306 1584 15312
rect 126 15272 138 15306
rect 1572 15272 1584 15306
rect 126 15266 900 15272
rect 894 15263 900 15266
rect 1548 15266 1584 15272
rect 1548 15263 1554 15266
rect 156 15226 162 15229
rect 126 15220 162 15226
rect 810 15226 816 15229
rect 810 15220 1584 15226
rect 126 15186 138 15220
rect 1572 15186 1584 15220
rect 126 15180 162 15186
rect 156 15177 162 15180
rect 810 15180 1584 15186
rect 810 15177 816 15180
rect 894 15140 900 15143
rect 126 15134 900 15140
rect 1548 15140 1554 15143
rect 1548 15134 1584 15140
rect 126 15100 138 15134
rect 1572 15100 1584 15134
rect 126 15094 900 15100
rect 894 15091 900 15094
rect 1548 15094 1584 15100
rect 1548 15091 1554 15094
rect 156 15054 162 15057
rect 126 15048 162 15054
rect 810 15054 816 15057
rect 810 15048 1584 15054
rect 126 15014 138 15048
rect 1572 15014 1584 15048
rect 126 15008 162 15014
rect 156 15005 162 15008
rect 810 15008 1584 15014
rect 810 15005 816 15008
rect 894 14968 900 14971
rect 126 14962 900 14968
rect 1548 14968 1554 14971
rect 1548 14962 1584 14968
rect 126 14928 138 14962
rect 1572 14928 1584 14962
rect 126 14922 900 14928
rect 894 14919 900 14922
rect 1548 14922 1584 14928
rect 1548 14919 1554 14922
rect 156 14882 162 14885
rect 126 14876 162 14882
rect 810 14882 816 14885
rect 810 14876 1584 14882
rect 126 14842 138 14876
rect 1572 14842 1584 14876
rect 126 14836 162 14842
rect 156 14833 162 14836
rect 810 14836 1584 14842
rect 810 14833 816 14836
rect 894 14796 900 14799
rect 126 14790 900 14796
rect 1548 14796 1554 14799
rect 1548 14790 1584 14796
rect 126 14756 138 14790
rect 1572 14756 1584 14790
rect 126 14750 900 14756
rect 894 14747 900 14750
rect 1548 14750 1584 14756
rect 1548 14747 1554 14750
rect 156 14710 162 14713
rect 126 14704 162 14710
rect 810 14710 816 14713
rect 810 14704 1584 14710
rect 126 14670 138 14704
rect 1572 14670 1584 14704
rect 126 14664 162 14670
rect 156 14661 162 14664
rect 810 14664 1584 14670
rect 810 14661 816 14664
rect 894 14624 900 14627
rect 126 14618 900 14624
rect 1548 14624 1554 14627
rect 1548 14618 1584 14624
rect 126 14584 138 14618
rect 1572 14584 1584 14618
rect 126 14578 900 14584
rect 894 14575 900 14578
rect 1548 14578 1584 14584
rect 1548 14575 1554 14578
rect 156 14538 162 14541
rect 126 14532 162 14538
rect 810 14538 816 14541
rect 810 14532 1584 14538
rect 126 14498 138 14532
rect 1572 14498 1584 14532
rect 126 14492 162 14498
rect 156 14489 162 14492
rect 810 14492 1584 14498
rect 810 14489 816 14492
rect 894 14452 900 14455
rect 126 14446 900 14452
rect 1548 14452 1554 14455
rect 1548 14446 1584 14452
rect 126 14412 138 14446
rect 1572 14412 1584 14446
rect 126 14406 900 14412
rect 894 14403 900 14406
rect 1548 14406 1584 14412
rect 1548 14403 1554 14406
rect 156 14366 162 14369
rect 126 14360 162 14366
rect 810 14366 816 14369
rect 810 14360 1584 14366
rect 126 14326 138 14360
rect 1572 14326 1584 14360
rect 126 14320 162 14326
rect 156 14317 162 14320
rect 810 14320 1584 14326
rect 810 14317 816 14320
rect 894 14280 900 14283
rect 126 14274 900 14280
rect 1548 14280 1554 14283
rect 1548 14274 1584 14280
rect 126 14240 138 14274
rect 1572 14240 1584 14274
rect 126 14234 900 14240
rect 894 14231 900 14234
rect 1548 14234 1584 14240
rect 1548 14231 1554 14234
rect 156 14194 162 14197
rect 126 14188 162 14194
rect 810 14194 816 14197
rect 810 14188 1584 14194
rect 126 14154 138 14188
rect 1572 14154 1584 14188
rect 126 14148 162 14154
rect 156 14145 162 14148
rect 810 14148 1584 14154
rect 810 14145 816 14148
rect 894 14108 900 14111
rect 126 14102 900 14108
rect 1548 14108 1554 14111
rect 1548 14102 1584 14108
rect 126 14068 138 14102
rect 1572 14068 1584 14102
rect 126 14062 900 14068
rect 894 14059 900 14062
rect 1548 14062 1584 14068
rect 1548 14059 1554 14062
rect 156 14022 162 14025
rect 126 14016 162 14022
rect 810 14022 816 14025
rect 810 14016 1584 14022
rect 126 13982 138 14016
rect 1572 13982 1584 14016
rect 126 13976 162 13982
rect 156 13973 162 13976
rect 810 13976 1584 13982
rect 810 13973 816 13976
rect 894 13936 900 13939
rect 126 13930 900 13936
rect 1548 13936 1554 13939
rect 1548 13930 1584 13936
rect 126 13896 138 13930
rect 1572 13896 1584 13930
rect 126 13890 900 13896
rect 894 13887 900 13890
rect 1548 13890 1584 13896
rect 1548 13887 1554 13890
rect 156 13850 162 13853
rect 126 13844 162 13850
rect 810 13850 816 13853
rect 810 13844 1584 13850
rect 126 13810 138 13844
rect 1572 13810 1584 13844
rect 126 13804 162 13810
rect 156 13801 162 13804
rect 810 13804 1584 13810
rect 810 13801 816 13804
rect 894 13764 900 13767
rect 126 13758 900 13764
rect 1548 13764 1554 13767
rect 1548 13758 1584 13764
rect 126 13724 138 13758
rect 1572 13724 1584 13758
rect 126 13718 900 13724
rect 894 13715 900 13718
rect 1548 13718 1584 13724
rect 1548 13715 1554 13718
rect 156 13678 162 13681
rect 126 13672 162 13678
rect 810 13678 816 13681
rect 810 13672 1584 13678
rect 126 13638 138 13672
rect 1572 13638 1584 13672
rect 126 13632 162 13638
rect 156 13629 162 13632
rect 810 13632 1584 13638
rect 810 13629 816 13632
rect 894 13592 900 13595
rect 126 13586 900 13592
rect 1548 13592 1554 13595
rect 1548 13586 1584 13592
rect 126 13552 138 13586
rect 1572 13552 1584 13586
rect 126 13546 900 13552
rect 894 13543 900 13546
rect 1548 13546 1584 13552
rect 1548 13543 1554 13546
rect 156 13506 162 13509
rect 126 13500 162 13506
rect 810 13506 816 13509
rect 810 13500 1584 13506
rect 126 13466 138 13500
rect 1572 13466 1584 13500
rect 126 13460 162 13466
rect 156 13457 162 13460
rect 810 13460 1584 13466
rect 810 13457 816 13460
rect 894 13420 900 13423
rect 126 13414 900 13420
rect 1548 13420 1554 13423
rect 1548 13414 1584 13420
rect 126 13380 138 13414
rect 1572 13380 1584 13414
rect 126 13374 900 13380
rect 894 13371 900 13374
rect 1548 13374 1584 13380
rect 1548 13371 1554 13374
rect 156 13334 162 13337
rect 126 13328 162 13334
rect 810 13334 816 13337
rect 810 13328 1584 13334
rect 126 13294 138 13328
rect 1572 13294 1584 13328
rect 126 13288 162 13294
rect 156 13285 162 13288
rect 810 13288 1584 13294
rect 810 13285 816 13288
rect 894 13248 900 13251
rect 126 13242 900 13248
rect 1548 13248 1554 13251
rect 1548 13242 1584 13248
rect 126 13208 138 13242
rect 1572 13208 1584 13242
rect 126 13202 900 13208
rect 894 13199 900 13202
rect 1548 13202 1584 13208
rect 1548 13199 1554 13202
rect 156 13162 162 13165
rect 126 13156 162 13162
rect 810 13162 816 13165
rect 810 13156 1584 13162
rect 126 13122 138 13156
rect 1572 13122 1584 13156
rect 126 13116 162 13122
rect 156 13113 162 13116
rect 810 13116 1584 13122
rect 810 13113 816 13116
rect 894 13076 900 13079
rect 126 13070 900 13076
rect 1548 13076 1554 13079
rect 1548 13070 1584 13076
rect 126 13036 138 13070
rect 1572 13036 1584 13070
rect 126 13030 900 13036
rect 894 13027 900 13030
rect 1548 13030 1584 13036
rect 1548 13027 1554 13030
rect 156 12990 162 12993
rect 126 12984 162 12990
rect 810 12990 816 12993
rect 810 12984 1584 12990
rect 126 12950 138 12984
rect 1572 12950 1584 12984
rect 126 12944 162 12950
rect 156 12941 162 12944
rect 810 12944 1584 12950
rect 810 12941 816 12944
rect 894 12904 900 12907
rect 126 12898 900 12904
rect 1548 12904 1554 12907
rect 1548 12898 1584 12904
rect 126 12864 138 12898
rect 1572 12864 1584 12898
rect 126 12858 900 12864
rect 894 12855 900 12858
rect 1548 12858 1584 12864
rect 1548 12855 1554 12858
rect 156 12818 162 12821
rect 126 12812 162 12818
rect 810 12818 816 12821
rect 810 12812 1584 12818
rect 126 12778 138 12812
rect 1572 12778 1584 12812
rect 126 12772 162 12778
rect 156 12769 162 12772
rect 810 12772 1584 12778
rect 810 12769 816 12772
rect 894 12732 900 12735
rect 126 12726 900 12732
rect 1548 12732 1554 12735
rect 1548 12726 1584 12732
rect 126 12692 138 12726
rect 1572 12692 1584 12726
rect 126 12686 900 12692
rect 894 12683 900 12686
rect 1548 12686 1584 12692
rect 1548 12683 1554 12686
rect 156 12646 162 12649
rect 126 12640 162 12646
rect 810 12646 816 12649
rect 810 12640 1584 12646
rect 126 12606 138 12640
rect 1572 12606 1584 12640
rect 126 12600 162 12606
rect 156 12597 162 12600
rect 810 12600 1584 12606
rect 810 12597 816 12600
rect 894 12560 900 12563
rect 126 12554 900 12560
rect 1548 12560 1554 12563
rect 1548 12554 1584 12560
rect 126 12520 138 12554
rect 1572 12520 1584 12554
rect 126 12514 900 12520
rect 894 12511 900 12514
rect 1548 12514 1584 12520
rect 1548 12511 1554 12514
rect 156 12474 162 12477
rect 126 12468 162 12474
rect 810 12474 816 12477
rect 810 12468 1584 12474
rect 126 12434 138 12468
rect 1572 12434 1584 12468
rect 126 12428 162 12434
rect 156 12425 162 12428
rect 810 12428 1584 12434
rect 810 12425 816 12428
rect 894 12388 900 12391
rect 126 12382 900 12388
rect 1548 12388 1554 12391
rect 1548 12382 1584 12388
rect 126 12348 138 12382
rect 1572 12348 1584 12382
rect 126 12342 900 12348
rect 894 12339 900 12342
rect 1548 12342 1584 12348
rect 1548 12339 1554 12342
rect 156 12302 162 12305
rect 126 12296 162 12302
rect 810 12302 816 12305
rect 810 12296 1584 12302
rect 126 12262 138 12296
rect 1572 12262 1584 12296
rect 126 12256 162 12262
rect 156 12253 162 12256
rect 810 12256 1584 12262
rect 810 12253 816 12256
rect 894 12216 900 12219
rect 126 12210 900 12216
rect 1548 12216 1554 12219
rect 1548 12210 1584 12216
rect 126 12176 138 12210
rect 1572 12176 1584 12210
rect 126 12170 900 12176
rect 894 12167 900 12170
rect 1548 12170 1584 12176
rect 1548 12167 1554 12170
rect 156 12130 162 12133
rect 126 12124 162 12130
rect 810 12130 816 12133
rect 810 12124 1584 12130
rect 126 12090 138 12124
rect 1572 12090 1584 12124
rect 126 12084 162 12090
rect 156 12081 162 12084
rect 810 12084 1584 12090
rect 810 12081 816 12084
rect 894 12044 900 12047
rect 126 12038 900 12044
rect 1548 12044 1554 12047
rect 1548 12038 1584 12044
rect 126 12004 138 12038
rect 1572 12004 1584 12038
rect 126 11998 900 12004
rect 894 11995 900 11998
rect 1548 11998 1584 12004
rect 1548 11995 1554 11998
rect 156 11958 162 11961
rect 126 11952 162 11958
rect 810 11958 816 11961
rect 810 11952 1584 11958
rect 126 11918 138 11952
rect 1572 11918 1584 11952
rect 126 11912 162 11918
rect 156 11909 162 11912
rect 810 11912 1584 11918
rect 810 11909 816 11912
rect 894 11872 900 11875
rect 126 11866 900 11872
rect 1548 11872 1554 11875
rect 1548 11866 1584 11872
rect 126 11832 138 11866
rect 1572 11832 1584 11866
rect 126 11826 900 11832
rect 894 11823 900 11826
rect 1548 11826 1584 11832
rect 1548 11823 1554 11826
rect 156 11786 162 11789
rect 126 11780 162 11786
rect 810 11786 816 11789
rect 810 11780 1584 11786
rect 126 11746 138 11780
rect 1572 11746 1584 11780
rect 126 11740 162 11746
rect 156 11737 162 11740
rect 810 11740 1584 11746
rect 810 11737 816 11740
rect 894 11700 900 11703
rect 126 11694 900 11700
rect 1548 11700 1554 11703
rect 1548 11694 1584 11700
rect 126 11660 138 11694
rect 1572 11660 1584 11694
rect 126 11654 900 11660
rect 894 11651 900 11654
rect 1548 11654 1584 11660
rect 1548 11651 1554 11654
rect 156 11614 162 11617
rect 126 11608 162 11614
rect 810 11614 816 11617
rect 810 11608 1584 11614
rect 126 11574 138 11608
rect 1572 11574 1584 11608
rect 126 11568 162 11574
rect 156 11565 162 11568
rect 810 11568 1584 11574
rect 810 11565 816 11568
rect 894 11528 900 11531
rect 126 11522 900 11528
rect 1548 11528 1554 11531
rect 1548 11522 1584 11528
rect 126 11488 138 11522
rect 1572 11488 1584 11522
rect 126 11482 900 11488
rect 894 11479 900 11482
rect 1548 11482 1584 11488
rect 1548 11479 1554 11482
rect 156 11442 162 11445
rect 126 11436 162 11442
rect 810 11442 816 11445
rect 810 11436 1584 11442
rect 126 11402 138 11436
rect 1572 11402 1584 11436
rect 126 11396 162 11402
rect 156 11393 162 11396
rect 810 11396 1584 11402
rect 810 11393 816 11396
rect 894 11356 900 11359
rect 126 11350 900 11356
rect 1548 11356 1554 11359
rect 1548 11350 1584 11356
rect 126 11316 138 11350
rect 1572 11316 1584 11350
rect 126 11310 900 11316
rect 894 11307 900 11310
rect 1548 11310 1584 11316
rect 1548 11307 1554 11310
rect 156 11270 162 11273
rect 126 11264 162 11270
rect 810 11270 816 11273
rect 810 11264 1584 11270
rect 126 11230 138 11264
rect 1572 11230 1584 11264
rect 126 11224 162 11230
rect 156 11221 162 11224
rect 810 11224 1584 11230
rect 810 11221 816 11224
rect 894 11184 900 11187
rect 126 11178 900 11184
rect 1548 11184 1554 11187
rect 1548 11178 1584 11184
rect 126 11144 138 11178
rect 1572 11144 1584 11178
rect 126 11138 900 11144
rect 894 11135 900 11138
rect 1548 11138 1584 11144
rect 1548 11135 1554 11138
rect 156 11098 162 11101
rect 126 11092 162 11098
rect 810 11098 816 11101
rect 810 11092 1584 11098
rect 126 11058 138 11092
rect 1572 11058 1584 11092
rect 126 11052 162 11058
rect 156 11049 162 11052
rect 810 11052 1584 11058
rect 810 11049 816 11052
rect 894 11012 900 11015
rect 126 11006 900 11012
rect 1548 11012 1554 11015
rect 1548 11006 1584 11012
rect 126 10972 138 11006
rect 1572 10972 1584 11006
rect 126 10966 900 10972
rect 894 10963 900 10966
rect 1548 10966 1584 10972
rect 1548 10963 1554 10966
rect 156 10926 162 10929
rect 126 10920 162 10926
rect 810 10926 816 10929
rect 810 10920 1584 10926
rect 126 10886 138 10920
rect 1572 10886 1584 10920
rect 126 10880 162 10886
rect 156 10877 162 10880
rect 810 10880 1584 10886
rect 810 10877 816 10880
rect 894 10840 900 10843
rect 126 10834 900 10840
rect 1548 10840 1554 10843
rect 1548 10834 1584 10840
rect 126 10800 138 10834
rect 1572 10800 1584 10834
rect 126 10794 900 10800
rect 894 10791 900 10794
rect 1548 10794 1584 10800
rect 1548 10791 1554 10794
rect 156 10754 162 10757
rect 126 10748 162 10754
rect 810 10754 816 10757
rect 810 10748 1584 10754
rect 126 10714 138 10748
rect 1572 10714 1584 10748
rect 126 10708 162 10714
rect 156 10705 162 10708
rect 810 10708 1584 10714
rect 810 10705 816 10708
rect 894 10668 900 10671
rect 126 10662 900 10668
rect 1548 10668 1554 10671
rect 1548 10662 1584 10668
rect 126 10628 138 10662
rect 1572 10628 1584 10662
rect 126 10622 900 10628
rect 894 10619 900 10622
rect 1548 10622 1584 10628
rect 1548 10619 1554 10622
rect 156 10582 162 10585
rect 126 10576 162 10582
rect 810 10582 816 10585
rect 810 10576 1584 10582
rect 126 10542 138 10576
rect 1572 10542 1584 10576
rect 126 10536 162 10542
rect 156 10533 162 10536
rect 810 10536 1584 10542
rect 810 10533 816 10536
rect 894 10496 900 10499
rect 126 10490 900 10496
rect 1548 10496 1554 10499
rect 1548 10490 1584 10496
rect 126 10456 138 10490
rect 1572 10456 1584 10490
rect 126 10450 900 10456
rect 894 10447 900 10450
rect 1548 10450 1584 10456
rect 1548 10447 1554 10450
rect 156 10410 162 10413
rect 126 10404 162 10410
rect 810 10410 816 10413
rect 810 10404 1584 10410
rect 126 10370 138 10404
rect 1572 10370 1584 10404
rect 126 10364 162 10370
rect 156 10361 162 10364
rect 810 10364 1584 10370
rect 810 10361 816 10364
rect 894 10324 900 10327
rect 126 10318 900 10324
rect 1548 10324 1554 10327
rect 1548 10318 1584 10324
rect 126 10284 138 10318
rect 1572 10284 1584 10318
rect 126 10278 900 10284
rect 894 10275 900 10278
rect 1548 10278 1584 10284
rect 1548 10275 1554 10278
rect 156 10238 162 10241
rect 126 10232 162 10238
rect 810 10238 816 10241
rect 810 10232 1584 10238
rect 126 10198 138 10232
rect 1572 10198 1584 10232
rect 126 10192 162 10198
rect 156 10189 162 10192
rect 810 10192 1584 10198
rect 810 10189 816 10192
rect 894 10152 900 10155
rect 126 10146 900 10152
rect 1548 10152 1554 10155
rect 1548 10146 1584 10152
rect 126 10112 138 10146
rect 1572 10112 1584 10146
rect 126 10106 900 10112
rect 894 10103 900 10106
rect 1548 10106 1584 10112
rect 1548 10103 1554 10106
rect 156 10066 162 10069
rect 126 10060 162 10066
rect 810 10066 816 10069
rect 810 10060 1584 10066
rect 126 10026 138 10060
rect 1572 10026 1584 10060
rect 126 10020 162 10026
rect 156 10017 162 10020
rect 810 10020 1584 10026
rect 810 10017 816 10020
rect 894 9980 900 9983
rect 126 9974 900 9980
rect 1548 9980 1554 9983
rect 1548 9974 1584 9980
rect 126 9940 138 9974
rect 1572 9940 1584 9974
rect 126 9934 900 9940
rect 894 9931 900 9934
rect 1548 9934 1584 9940
rect 1548 9931 1554 9934
rect 156 9894 162 9897
rect 126 9888 162 9894
rect 810 9894 816 9897
rect 810 9888 1584 9894
rect 126 9854 138 9888
rect 1572 9854 1584 9888
rect 126 9848 162 9854
rect 156 9845 162 9848
rect 810 9848 1584 9854
rect 810 9845 816 9848
rect 894 9808 900 9811
rect 126 9802 900 9808
rect 1548 9808 1554 9811
rect 1548 9802 1584 9808
rect 126 9768 138 9802
rect 1572 9768 1584 9802
rect 126 9762 900 9768
rect 894 9759 900 9762
rect 1548 9762 1584 9768
rect 1548 9759 1554 9762
rect 156 9722 162 9725
rect 126 9716 162 9722
rect 810 9722 816 9725
rect 810 9716 1584 9722
rect 126 9682 138 9716
rect 1572 9682 1584 9716
rect 126 9676 162 9682
rect 156 9673 162 9676
rect 810 9676 1584 9682
rect 810 9673 816 9676
rect 894 9636 900 9639
rect 126 9630 900 9636
rect 1548 9636 1554 9639
rect 1548 9630 1584 9636
rect 126 9596 138 9630
rect 1572 9596 1584 9630
rect 126 9590 900 9596
rect 894 9587 900 9590
rect 1548 9590 1584 9596
rect 1548 9587 1554 9590
rect 156 9550 162 9553
rect 126 9544 162 9550
rect 810 9550 816 9553
rect 810 9544 1584 9550
rect 126 9510 138 9544
rect 1572 9510 1584 9544
rect 126 9504 162 9510
rect 156 9501 162 9504
rect 810 9504 1584 9510
rect 810 9501 816 9504
rect 894 9464 900 9467
rect 126 9458 900 9464
rect 1548 9464 1554 9467
rect 1548 9458 1584 9464
rect 126 9424 138 9458
rect 1572 9424 1584 9458
rect 126 9418 900 9424
rect 894 9415 900 9418
rect 1548 9418 1584 9424
rect 1548 9415 1554 9418
rect 156 9378 162 9381
rect 126 9372 162 9378
rect 810 9378 816 9381
rect 810 9372 1584 9378
rect 126 9338 138 9372
rect 1572 9338 1584 9372
rect 126 9332 162 9338
rect 156 9329 162 9332
rect 810 9332 1584 9338
rect 810 9329 816 9332
rect 894 9292 900 9295
rect 126 9286 900 9292
rect 1548 9292 1554 9295
rect 1548 9286 1584 9292
rect 126 9252 138 9286
rect 1572 9252 1584 9286
rect 126 9246 900 9252
rect 894 9243 900 9246
rect 1548 9246 1584 9252
rect 1548 9243 1554 9246
rect 156 9206 162 9209
rect 126 9200 162 9206
rect 810 9206 816 9209
rect 810 9200 1584 9206
rect 126 9166 138 9200
rect 1572 9166 1584 9200
rect 126 9160 162 9166
rect 156 9157 162 9160
rect 810 9160 1584 9166
rect 810 9157 816 9160
rect 894 9120 900 9123
rect 126 9114 900 9120
rect 1548 9120 1554 9123
rect 1548 9114 1584 9120
rect 126 9080 138 9114
rect 1572 9080 1584 9114
rect 126 9074 900 9080
rect 894 9071 900 9074
rect 1548 9074 1584 9080
rect 1548 9071 1554 9074
rect 156 9034 162 9037
rect 126 9028 162 9034
rect 810 9034 816 9037
rect 810 9028 1584 9034
rect 126 8994 138 9028
rect 1572 8994 1584 9028
rect 126 8988 162 8994
rect 156 8985 162 8988
rect 810 8988 1584 8994
rect 810 8985 816 8988
rect 894 8948 900 8951
rect 126 8942 900 8948
rect 1548 8948 1554 8951
rect 1548 8942 1584 8948
rect 126 8908 138 8942
rect 1572 8908 1584 8942
rect 126 8902 900 8908
rect 894 8899 900 8902
rect 1548 8902 1584 8908
rect 1548 8899 1554 8902
rect 156 8862 162 8865
rect 126 8856 162 8862
rect 810 8862 816 8865
rect 810 8856 1584 8862
rect 126 8822 138 8856
rect 1572 8822 1584 8856
rect 126 8816 162 8822
rect 156 8813 162 8816
rect 810 8816 1584 8822
rect 810 8813 816 8816
rect 894 8776 900 8779
rect 126 8770 900 8776
rect 1548 8776 1554 8779
rect 1548 8770 1584 8776
rect 126 8736 138 8770
rect 1572 8736 1584 8770
rect 126 8730 900 8736
rect 894 8727 900 8730
rect 1548 8730 1584 8736
rect 1548 8727 1554 8730
rect 156 8690 162 8693
rect 126 8684 162 8690
rect 810 8690 816 8693
rect 810 8684 1584 8690
rect 126 8650 138 8684
rect 1572 8650 1584 8684
rect 126 8644 162 8650
rect 156 8641 162 8644
rect 810 8644 1584 8650
rect 810 8641 816 8644
rect 894 8604 900 8607
rect 126 8598 900 8604
rect 1548 8604 1554 8607
rect 1548 8598 1584 8604
rect 126 8564 138 8598
rect 1572 8564 1584 8598
rect 126 8558 900 8564
rect 894 8555 900 8558
rect 1548 8558 1584 8564
rect 1548 8555 1554 8558
rect 156 8518 162 8521
rect 126 8512 162 8518
rect 810 8518 816 8521
rect 810 8512 1584 8518
rect 126 8478 138 8512
rect 1572 8478 1584 8512
rect 126 8472 162 8478
rect 156 8469 162 8472
rect 810 8472 1584 8478
rect 810 8469 816 8472
rect 894 8432 900 8435
rect 126 8426 900 8432
rect 1548 8432 1554 8435
rect 1548 8426 1584 8432
rect 126 8392 138 8426
rect 1572 8392 1584 8426
rect 126 8386 900 8392
rect 894 8383 900 8386
rect 1548 8386 1584 8392
rect 1548 8383 1554 8386
rect 156 8346 162 8349
rect 126 8340 162 8346
rect 810 8346 816 8349
rect 810 8340 1584 8346
rect 126 8306 138 8340
rect 1572 8306 1584 8340
rect 126 8300 162 8306
rect 156 8297 162 8300
rect 810 8300 1584 8306
rect 810 8297 816 8300
rect 894 8260 900 8263
rect 126 8254 900 8260
rect 1548 8260 1554 8263
rect 1548 8254 1584 8260
rect 126 8220 138 8254
rect 1572 8220 1584 8254
rect 126 8214 900 8220
rect 894 8211 900 8214
rect 1548 8214 1584 8220
rect 1548 8211 1554 8214
rect 156 8174 162 8177
rect 126 8168 162 8174
rect 810 8174 816 8177
rect 810 8168 1584 8174
rect 126 8134 138 8168
rect 1572 8134 1584 8168
rect 126 8128 162 8134
rect 156 8125 162 8128
rect 810 8128 1584 8134
rect 810 8125 816 8128
rect 894 8088 900 8091
rect 126 8082 900 8088
rect 1548 8088 1554 8091
rect 1548 8082 1584 8088
rect 126 8048 138 8082
rect 1572 8048 1584 8082
rect 126 8042 900 8048
rect 894 8039 900 8042
rect 1548 8042 1584 8048
rect 1548 8039 1554 8042
rect 156 8002 162 8005
rect 126 7996 162 8002
rect 810 8002 816 8005
rect 810 7996 1584 8002
rect 126 7962 138 7996
rect 1572 7962 1584 7996
rect 126 7956 162 7962
rect 156 7953 162 7956
rect 810 7956 1584 7962
rect 810 7953 816 7956
rect 894 7916 900 7919
rect 126 7910 900 7916
rect 1548 7916 1554 7919
rect 1548 7910 1584 7916
rect 126 7876 138 7910
rect 1572 7876 1584 7910
rect 126 7870 900 7876
rect 894 7867 900 7870
rect 1548 7870 1584 7876
rect 1548 7867 1554 7870
rect 156 7830 162 7833
rect 126 7824 162 7830
rect 810 7830 816 7833
rect 810 7824 1584 7830
rect 126 7790 138 7824
rect 1572 7790 1584 7824
rect 126 7784 162 7790
rect 156 7781 162 7784
rect 810 7784 1584 7790
rect 810 7781 816 7784
rect 894 7744 900 7747
rect 126 7738 900 7744
rect 1548 7744 1554 7747
rect 1548 7738 1584 7744
rect 126 7704 138 7738
rect 1572 7704 1584 7738
rect 126 7698 900 7704
rect 894 7695 900 7698
rect 1548 7698 1584 7704
rect 1548 7695 1554 7698
rect 156 7658 162 7661
rect 126 7652 162 7658
rect 810 7658 816 7661
rect 810 7652 1584 7658
rect 126 7618 138 7652
rect 1572 7618 1584 7652
rect 126 7612 162 7618
rect 156 7609 162 7612
rect 810 7612 1584 7618
rect 810 7609 816 7612
rect 894 7572 900 7575
rect 126 7566 900 7572
rect 1548 7572 1554 7575
rect 1548 7566 1584 7572
rect 126 7532 138 7566
rect 1572 7532 1584 7566
rect 126 7526 900 7532
rect 894 7523 900 7526
rect 1548 7526 1584 7532
rect 1548 7523 1554 7526
rect 156 7486 162 7489
rect 126 7480 162 7486
rect 810 7486 816 7489
rect 810 7480 1584 7486
rect 126 7446 138 7480
rect 1572 7446 1584 7480
rect 126 7440 162 7446
rect 156 7437 162 7440
rect 810 7440 1584 7446
rect 810 7437 816 7440
rect 894 7400 900 7403
rect 126 7394 900 7400
rect 1548 7400 1554 7403
rect 1548 7394 1584 7400
rect 126 7360 138 7394
rect 1572 7360 1584 7394
rect 126 7354 900 7360
rect 894 7351 900 7354
rect 1548 7354 1584 7360
rect 1548 7351 1554 7354
rect 156 7314 162 7317
rect 126 7308 162 7314
rect 810 7314 816 7317
rect 810 7308 1584 7314
rect 126 7274 138 7308
rect 1572 7274 1584 7308
rect 126 7268 162 7274
rect 156 7265 162 7268
rect 810 7268 1584 7274
rect 810 7265 816 7268
rect 894 7228 900 7231
rect 126 7222 900 7228
rect 1548 7228 1554 7231
rect 1548 7222 1584 7228
rect 126 7188 138 7222
rect 1572 7188 1584 7222
rect 126 7182 900 7188
rect 894 7179 900 7182
rect 1548 7182 1584 7188
rect 1548 7179 1554 7182
rect 156 7142 162 7145
rect 126 7136 162 7142
rect 810 7142 816 7145
rect 810 7136 1584 7142
rect 126 7102 138 7136
rect 1572 7102 1584 7136
rect 126 7096 162 7102
rect 156 7093 162 7096
rect 810 7096 1584 7102
rect 810 7093 816 7096
rect 894 7056 900 7059
rect 126 7050 900 7056
rect 1548 7056 1554 7059
rect 1548 7050 1584 7056
rect 126 7016 138 7050
rect 1572 7016 1584 7050
rect 126 7010 900 7016
rect 894 7007 900 7010
rect 1548 7010 1584 7016
rect 1548 7007 1554 7010
rect 156 6970 162 6973
rect 126 6964 162 6970
rect 810 6970 816 6973
rect 810 6964 1584 6970
rect 126 6930 138 6964
rect 1572 6930 1584 6964
rect 126 6924 162 6930
rect 156 6921 162 6924
rect 810 6924 1584 6930
rect 810 6921 816 6924
rect 894 6884 900 6887
rect 126 6878 900 6884
rect 1548 6884 1554 6887
rect 1548 6878 1584 6884
rect 126 6844 138 6878
rect 1572 6844 1584 6878
rect 126 6838 900 6844
rect 894 6835 900 6838
rect 1548 6838 1584 6844
rect 1548 6835 1554 6838
rect 156 6798 162 6801
rect 126 6792 162 6798
rect 810 6798 816 6801
rect 810 6792 1584 6798
rect 126 6758 138 6792
rect 1572 6758 1584 6792
rect 126 6752 162 6758
rect 156 6749 162 6752
rect 810 6752 1584 6758
rect 810 6749 816 6752
rect 894 6712 900 6715
rect 126 6706 900 6712
rect 1548 6712 1554 6715
rect 1548 6706 1584 6712
rect 126 6672 138 6706
rect 1572 6672 1584 6706
rect 126 6666 900 6672
rect 894 6663 900 6666
rect 1548 6666 1584 6672
rect 1548 6663 1554 6666
rect 156 6626 162 6629
rect 126 6620 162 6626
rect 810 6626 816 6629
rect 810 6620 1584 6626
rect 126 6586 138 6620
rect 1572 6586 1584 6620
rect 126 6580 162 6586
rect 156 6577 162 6580
rect 810 6580 1584 6586
rect 810 6577 816 6580
rect 894 6540 900 6543
rect 126 6534 900 6540
rect 1548 6540 1554 6543
rect 1548 6534 1584 6540
rect 126 6500 138 6534
rect 1572 6500 1584 6534
rect 126 6494 900 6500
rect 894 6491 900 6494
rect 1548 6494 1584 6500
rect 1548 6491 1554 6494
rect 156 6454 162 6457
rect 126 6448 162 6454
rect 810 6454 816 6457
rect 810 6448 1584 6454
rect 126 6414 138 6448
rect 1572 6414 1584 6448
rect 126 6408 162 6414
rect 156 6405 162 6408
rect 810 6408 1584 6414
rect 810 6405 816 6408
rect 894 6368 900 6371
rect 126 6362 900 6368
rect 1548 6368 1554 6371
rect 1548 6362 1584 6368
rect 126 6328 138 6362
rect 1572 6328 1584 6362
rect 126 6322 900 6328
rect 894 6319 900 6322
rect 1548 6322 1584 6328
rect 1548 6319 1554 6322
rect 156 6282 162 6285
rect 126 6276 162 6282
rect 810 6282 816 6285
rect 810 6276 1584 6282
rect 126 6242 138 6276
rect 1572 6242 1584 6276
rect 126 6236 162 6242
rect 156 6233 162 6236
rect 810 6236 1584 6242
rect 810 6233 816 6236
rect 894 6196 900 6199
rect 126 6190 900 6196
rect 1548 6196 1554 6199
rect 1548 6190 1584 6196
rect 126 6156 138 6190
rect 1572 6156 1584 6190
rect 126 6150 900 6156
rect 894 6147 900 6150
rect 1548 6150 1584 6156
rect 1548 6147 1554 6150
rect 156 6110 162 6113
rect 126 6104 162 6110
rect 810 6110 816 6113
rect 810 6104 1584 6110
rect 126 6070 138 6104
rect 1572 6070 1584 6104
rect 126 6064 162 6070
rect 156 6061 162 6064
rect 810 6064 1584 6070
rect 810 6061 816 6064
rect 894 6024 900 6027
rect 126 6018 900 6024
rect 1548 6024 1554 6027
rect 1548 6018 1584 6024
rect 126 5984 138 6018
rect 1572 5984 1584 6018
rect 126 5978 900 5984
rect 894 5975 900 5978
rect 1548 5978 1584 5984
rect 1548 5975 1554 5978
rect 156 5938 162 5941
rect 126 5932 162 5938
rect 810 5938 816 5941
rect 810 5932 1584 5938
rect 126 5898 138 5932
rect 1572 5898 1584 5932
rect 126 5892 162 5898
rect 156 5889 162 5892
rect 810 5892 1584 5898
rect 810 5889 816 5892
rect 894 5852 900 5855
rect 126 5846 900 5852
rect 1548 5852 1554 5855
rect 1548 5846 1584 5852
rect 126 5812 138 5846
rect 1572 5812 1584 5846
rect 126 5806 900 5812
rect 894 5803 900 5806
rect 1548 5806 1584 5812
rect 1548 5803 1554 5806
rect 156 5766 162 5769
rect 126 5760 162 5766
rect 810 5766 816 5769
rect 810 5760 1584 5766
rect 126 5726 138 5760
rect 1572 5726 1584 5760
rect 126 5720 162 5726
rect 156 5717 162 5720
rect 810 5720 1584 5726
rect 810 5717 816 5720
rect 894 5680 900 5683
rect 126 5674 900 5680
rect 1548 5680 1554 5683
rect 1548 5674 1584 5680
rect 126 5640 138 5674
rect 1572 5640 1584 5674
rect 126 5634 900 5640
rect 894 5631 900 5634
rect 1548 5634 1584 5640
rect 1548 5631 1554 5634
rect 156 5594 162 5597
rect 126 5588 162 5594
rect 810 5594 816 5597
rect 810 5588 1584 5594
rect 126 5554 138 5588
rect 1572 5554 1584 5588
rect 126 5548 162 5554
rect 156 5545 162 5548
rect 810 5548 1584 5554
rect 810 5545 816 5548
rect 894 5508 900 5511
rect 126 5502 900 5508
rect 1548 5508 1554 5511
rect 1548 5502 1584 5508
rect 126 5468 138 5502
rect 1572 5468 1584 5502
rect 126 5462 900 5468
rect 894 5459 900 5462
rect 1548 5462 1584 5468
rect 1548 5459 1554 5462
rect 156 5422 162 5425
rect 126 5416 162 5422
rect 810 5422 816 5425
rect 810 5416 1584 5422
rect 126 5382 138 5416
rect 1572 5382 1584 5416
rect 126 5376 162 5382
rect 156 5373 162 5376
rect 810 5376 1584 5382
rect 810 5373 816 5376
rect 894 5336 900 5339
rect 126 5330 900 5336
rect 1548 5336 1554 5339
rect 1548 5330 1584 5336
rect 126 5296 138 5330
rect 1572 5296 1584 5330
rect 126 5290 900 5296
rect 894 5287 900 5290
rect 1548 5290 1584 5296
rect 1548 5287 1554 5290
rect 156 5250 162 5253
rect 126 5244 162 5250
rect 810 5250 816 5253
rect 810 5244 1584 5250
rect 126 5210 138 5244
rect 1572 5210 1584 5244
rect 126 5204 162 5210
rect 156 5201 162 5204
rect 810 5204 1584 5210
rect 810 5201 816 5204
rect 894 5164 900 5167
rect 126 5158 900 5164
rect 1548 5164 1554 5167
rect 1548 5158 1584 5164
rect 126 5124 138 5158
rect 1572 5124 1584 5158
rect 126 5118 900 5124
rect 894 5115 900 5118
rect 1548 5118 1584 5124
rect 1548 5115 1554 5118
rect 156 5078 162 5081
rect 126 5072 162 5078
rect 810 5078 816 5081
rect 810 5072 1584 5078
rect 126 5038 138 5072
rect 1572 5038 1584 5072
rect 126 5032 162 5038
rect 156 5029 162 5032
rect 810 5032 1584 5038
rect 810 5029 816 5032
rect 894 4992 900 4995
rect 126 4986 900 4992
rect 1548 4992 1554 4995
rect 1548 4986 1584 4992
rect 126 4952 138 4986
rect 1572 4952 1584 4986
rect 126 4946 900 4952
rect 894 4943 900 4946
rect 1548 4946 1584 4952
rect 1548 4943 1554 4946
rect 156 4906 162 4909
rect 126 4900 162 4906
rect 810 4906 816 4909
rect 810 4900 1584 4906
rect 126 4866 138 4900
rect 1572 4866 1584 4900
rect 126 4860 162 4866
rect 156 4857 162 4860
rect 810 4860 1584 4866
rect 810 4857 816 4860
rect 894 4820 900 4823
rect 126 4814 900 4820
rect 1548 4820 1554 4823
rect 1548 4814 1584 4820
rect 126 4780 138 4814
rect 1572 4780 1584 4814
rect 126 4774 900 4780
rect 894 4771 900 4774
rect 1548 4774 1584 4780
rect 1548 4771 1554 4774
rect 156 4734 162 4737
rect 126 4728 162 4734
rect 810 4734 816 4737
rect 810 4728 1584 4734
rect 126 4694 138 4728
rect 1572 4694 1584 4728
rect 126 4688 162 4694
rect 156 4685 162 4688
rect 810 4688 1584 4694
rect 810 4685 816 4688
rect 894 4648 900 4651
rect 126 4642 900 4648
rect 1548 4648 1554 4651
rect 1548 4642 1584 4648
rect 126 4608 138 4642
rect 1572 4608 1584 4642
rect 126 4602 900 4608
rect 894 4599 900 4602
rect 1548 4602 1584 4608
rect 1548 4599 1554 4602
rect 156 4562 162 4565
rect 126 4556 162 4562
rect 810 4562 816 4565
rect 810 4556 1584 4562
rect 126 4522 138 4556
rect 1572 4522 1584 4556
rect 126 4516 162 4522
rect 156 4513 162 4516
rect 810 4516 1584 4522
rect 810 4513 816 4516
rect 894 4476 900 4479
rect 126 4470 900 4476
rect 1548 4476 1554 4479
rect 1548 4470 1584 4476
rect 126 4436 138 4470
rect 1572 4436 1584 4470
rect 126 4430 900 4436
rect 894 4427 900 4430
rect 1548 4430 1584 4436
rect 1548 4427 1554 4430
rect 156 4390 162 4393
rect 126 4384 162 4390
rect 810 4390 816 4393
rect 810 4384 1584 4390
rect 126 4350 138 4384
rect 1572 4350 1584 4384
rect 126 4344 162 4350
rect 156 4341 162 4344
rect 810 4344 1584 4350
rect 810 4341 816 4344
rect 894 4304 900 4307
rect 126 4298 900 4304
rect 1548 4304 1554 4307
rect 1548 4298 1584 4304
rect 126 4264 138 4298
rect 1572 4264 1584 4298
rect 126 4258 900 4264
rect 894 4255 900 4258
rect 1548 4258 1584 4264
rect 1548 4255 1554 4258
rect 156 4218 162 4221
rect 126 4212 162 4218
rect 810 4218 816 4221
rect 810 4212 1584 4218
rect 126 4178 138 4212
rect 1572 4178 1584 4212
rect 126 4172 162 4178
rect 156 4169 162 4172
rect 810 4172 1584 4178
rect 810 4169 816 4172
rect 894 4132 900 4135
rect 126 4126 900 4132
rect 1548 4132 1554 4135
rect 1548 4126 1584 4132
rect 126 4092 138 4126
rect 1572 4092 1584 4126
rect 126 4086 900 4092
rect 894 4083 900 4086
rect 1548 4086 1584 4092
rect 1548 4083 1554 4086
rect 156 4046 162 4049
rect 126 4040 162 4046
rect 810 4046 816 4049
rect 810 4040 1584 4046
rect 126 4006 138 4040
rect 1572 4006 1584 4040
rect 126 4000 162 4006
rect 156 3997 162 4000
rect 810 4000 1584 4006
rect 810 3997 816 4000
rect 894 3960 900 3963
rect 126 3954 900 3960
rect 1548 3960 1554 3963
rect 1548 3954 1584 3960
rect 126 3920 138 3954
rect 1572 3920 1584 3954
rect 126 3914 900 3920
rect 894 3911 900 3914
rect 1548 3914 1584 3920
rect 1548 3911 1554 3914
rect 156 3874 162 3877
rect 126 3868 162 3874
rect 810 3874 816 3877
rect 810 3868 1584 3874
rect 126 3834 138 3868
rect 1572 3834 1584 3868
rect 126 3828 162 3834
rect 156 3825 162 3828
rect 810 3828 1584 3834
rect 810 3825 816 3828
rect 894 3788 900 3791
rect 126 3782 900 3788
rect 1548 3788 1554 3791
rect 1548 3782 1584 3788
rect 126 3748 138 3782
rect 1572 3748 1584 3782
rect 126 3742 900 3748
rect 894 3739 900 3742
rect 1548 3742 1584 3748
rect 1548 3739 1554 3742
rect 156 3702 162 3705
rect 126 3696 162 3702
rect 810 3702 816 3705
rect 810 3696 1584 3702
rect 126 3662 138 3696
rect 1572 3662 1584 3696
rect 126 3656 162 3662
rect 156 3653 162 3656
rect 810 3656 1584 3662
rect 810 3653 816 3656
rect 894 3616 900 3619
rect 126 3610 900 3616
rect 1548 3616 1554 3619
rect 1548 3610 1584 3616
rect 126 3576 138 3610
rect 1572 3576 1584 3610
rect 126 3570 900 3576
rect 894 3567 900 3570
rect 1548 3570 1584 3576
rect 1548 3567 1554 3570
rect 156 3530 162 3533
rect 126 3524 162 3530
rect 810 3530 816 3533
rect 810 3524 1584 3530
rect 126 3490 138 3524
rect 1572 3490 1584 3524
rect 126 3484 162 3490
rect 156 3481 162 3484
rect 810 3484 1584 3490
rect 810 3481 816 3484
rect 894 3444 900 3447
rect 126 3438 900 3444
rect 1548 3444 1554 3447
rect 1548 3438 1584 3444
rect 126 3404 138 3438
rect 1572 3404 1584 3438
rect 126 3398 900 3404
rect 894 3395 900 3398
rect 1548 3398 1584 3404
rect 1548 3395 1554 3398
rect 156 3358 162 3361
rect 126 3352 162 3358
rect 810 3358 816 3361
rect 810 3352 1584 3358
rect 126 3318 138 3352
rect 1572 3318 1584 3352
rect 126 3312 162 3318
rect 156 3309 162 3312
rect 810 3312 1584 3318
rect 810 3309 816 3312
rect 894 3272 900 3275
rect 126 3266 900 3272
rect 1548 3272 1554 3275
rect 1548 3266 1584 3272
rect 126 3232 138 3266
rect 1572 3232 1584 3266
rect 126 3226 900 3232
rect 894 3223 900 3226
rect 1548 3226 1584 3232
rect 1548 3223 1554 3226
rect 156 3186 162 3189
rect 126 3180 162 3186
rect 810 3186 816 3189
rect 810 3180 1584 3186
rect 126 3146 138 3180
rect 1572 3146 1584 3180
rect 126 3140 162 3146
rect 156 3137 162 3140
rect 810 3140 1584 3146
rect 810 3137 816 3140
rect 894 3100 900 3103
rect 126 3094 900 3100
rect 1548 3100 1554 3103
rect 1548 3094 1584 3100
rect 126 3060 138 3094
rect 1572 3060 1584 3094
rect 126 3054 900 3060
rect 894 3051 900 3054
rect 1548 3054 1584 3060
rect 1548 3051 1554 3054
rect 156 3014 162 3017
rect 126 3008 162 3014
rect 810 3014 816 3017
rect 810 3008 1584 3014
rect 126 2974 138 3008
rect 1572 2974 1584 3008
rect 126 2968 162 2974
rect 156 2965 162 2968
rect 810 2968 1584 2974
rect 810 2965 816 2968
rect 894 2928 900 2931
rect 126 2922 900 2928
rect 1548 2928 1554 2931
rect 1548 2922 1584 2928
rect 126 2888 138 2922
rect 1572 2888 1584 2922
rect 126 2882 900 2888
rect 894 2879 900 2882
rect 1548 2882 1584 2888
rect 1548 2879 1554 2882
rect 156 2842 162 2845
rect 126 2836 162 2842
rect 810 2842 816 2845
rect 810 2836 1584 2842
rect 126 2802 138 2836
rect 1572 2802 1584 2836
rect 126 2796 162 2802
rect 156 2793 162 2796
rect 810 2796 1584 2802
rect 810 2793 816 2796
rect 894 2756 900 2759
rect 126 2750 900 2756
rect 1548 2756 1554 2759
rect 1548 2750 1584 2756
rect 126 2716 138 2750
rect 1572 2716 1584 2750
rect 126 2710 900 2716
rect 894 2707 900 2710
rect 1548 2710 1584 2716
rect 1548 2707 1554 2710
rect 156 2670 162 2673
rect 126 2664 162 2670
rect 810 2670 816 2673
rect 810 2664 1584 2670
rect 126 2630 138 2664
rect 1572 2630 1584 2664
rect 126 2624 162 2630
rect 156 2621 162 2624
rect 810 2624 1584 2630
rect 810 2621 816 2624
rect 894 2584 900 2587
rect 126 2578 900 2584
rect 1548 2584 1554 2587
rect 1548 2578 1584 2584
rect 126 2544 138 2578
rect 1572 2544 1584 2578
rect 126 2538 900 2544
rect 894 2535 900 2538
rect 1548 2538 1584 2544
rect 1548 2535 1554 2538
rect 156 2498 162 2501
rect 126 2492 162 2498
rect 810 2498 816 2501
rect 810 2492 1584 2498
rect 126 2458 138 2492
rect 1572 2458 1584 2492
rect 126 2452 162 2458
rect 156 2449 162 2452
rect 810 2452 1584 2458
rect 810 2449 816 2452
rect 894 2412 900 2415
rect 126 2406 900 2412
rect 1548 2412 1554 2415
rect 1548 2406 1584 2412
rect 126 2372 138 2406
rect 1572 2372 1584 2406
rect 126 2366 900 2372
rect 894 2363 900 2366
rect 1548 2366 1584 2372
rect 1548 2363 1554 2366
rect 156 2326 162 2329
rect 126 2320 162 2326
rect 810 2326 816 2329
rect 810 2320 1584 2326
rect 126 2286 138 2320
rect 1572 2286 1584 2320
rect 126 2280 162 2286
rect 156 2277 162 2280
rect 810 2280 1584 2286
rect 810 2277 816 2280
rect 894 2240 900 2243
rect 126 2234 900 2240
rect 1548 2240 1554 2243
rect 1548 2234 1584 2240
rect 126 2200 138 2234
rect 1572 2200 1584 2234
rect 126 2194 900 2200
rect 894 2191 900 2194
rect 1548 2194 1584 2200
rect 1548 2191 1554 2194
rect 156 2154 162 2157
rect 126 2148 162 2154
rect 810 2154 816 2157
rect 810 2148 1584 2154
rect 126 2114 138 2148
rect 1572 2114 1584 2148
rect 126 2108 162 2114
rect 156 2105 162 2108
rect 810 2108 1584 2114
rect 810 2105 816 2108
rect 894 2068 900 2071
rect 126 2062 900 2068
rect 1548 2068 1554 2071
rect 1548 2062 1584 2068
rect 126 2028 138 2062
rect 1572 2028 1584 2062
rect 126 2022 900 2028
rect 894 2019 900 2022
rect 1548 2022 1584 2028
rect 1548 2019 1554 2022
rect 156 1982 162 1985
rect 126 1976 162 1982
rect 810 1982 816 1985
rect 810 1976 1584 1982
rect 126 1942 138 1976
rect 1572 1942 1584 1976
rect 126 1936 162 1942
rect 156 1933 162 1936
rect 810 1936 1584 1942
rect 810 1933 816 1936
rect 894 1896 900 1899
rect 126 1890 900 1896
rect 1548 1896 1554 1899
rect 1548 1890 1584 1896
rect 126 1856 138 1890
rect 1572 1856 1584 1890
rect 126 1850 900 1856
rect 894 1847 900 1850
rect 1548 1850 1584 1856
rect 1548 1847 1554 1850
rect 156 1810 162 1813
rect 126 1804 162 1810
rect 810 1810 816 1813
rect 810 1804 1584 1810
rect 126 1770 138 1804
rect 1572 1770 1584 1804
rect 126 1764 162 1770
rect 156 1761 162 1764
rect 810 1764 1584 1770
rect 810 1761 816 1764
rect 894 1724 900 1727
rect 126 1718 900 1724
rect 1548 1724 1554 1727
rect 1548 1718 1584 1724
rect 126 1684 138 1718
rect 1572 1684 1584 1718
rect 126 1678 900 1684
rect 894 1675 900 1678
rect 1548 1678 1584 1684
rect 1548 1675 1554 1678
rect 156 1638 162 1641
rect 126 1632 162 1638
rect 810 1638 816 1641
rect 810 1632 1584 1638
rect 126 1598 138 1632
rect 1572 1598 1584 1632
rect 126 1592 162 1598
rect 156 1589 162 1592
rect 810 1592 1584 1598
rect 810 1589 816 1592
rect 894 1552 900 1555
rect 126 1546 900 1552
rect 1548 1552 1554 1555
rect 1548 1546 1584 1552
rect 126 1512 138 1546
rect 1572 1512 1584 1546
rect 126 1506 900 1512
rect 894 1503 900 1506
rect 1548 1506 1584 1512
rect 1548 1503 1554 1506
rect 156 1466 162 1469
rect 126 1460 162 1466
rect 810 1466 816 1469
rect 810 1460 1584 1466
rect 126 1426 138 1460
rect 1572 1426 1584 1460
rect 126 1420 162 1426
rect 156 1417 162 1420
rect 810 1420 1584 1426
rect 810 1417 816 1420
rect 894 1380 900 1383
rect 126 1374 900 1380
rect 1548 1380 1554 1383
rect 1548 1374 1584 1380
rect 126 1340 138 1374
rect 1572 1340 1584 1374
rect 126 1334 900 1340
rect 894 1331 900 1334
rect 1548 1334 1584 1340
rect 1548 1331 1554 1334
rect 156 1294 162 1297
rect 126 1288 162 1294
rect 810 1294 816 1297
rect 810 1288 1584 1294
rect 126 1254 138 1288
rect 1572 1254 1584 1288
rect 126 1248 162 1254
rect 156 1245 162 1248
rect 810 1248 1584 1254
rect 810 1245 816 1248
rect 894 1208 900 1211
rect 126 1202 900 1208
rect 1548 1208 1554 1211
rect 1548 1202 1584 1208
rect 126 1168 138 1202
rect 1572 1168 1584 1202
rect 126 1162 900 1168
rect 894 1159 900 1162
rect 1548 1162 1584 1168
rect 1548 1159 1554 1162
rect 156 1122 162 1125
rect 126 1116 162 1122
rect 810 1122 816 1125
rect 810 1116 1584 1122
rect 126 1082 138 1116
rect 1572 1082 1584 1116
rect 126 1076 162 1082
rect 156 1073 162 1076
rect 810 1076 1584 1082
rect 810 1073 816 1076
rect 894 1036 900 1039
rect 126 1030 900 1036
rect 1548 1036 1554 1039
rect 1548 1030 1584 1036
rect 126 996 138 1030
rect 1572 996 1584 1030
rect 126 990 900 996
rect 894 987 900 990
rect 1548 990 1584 996
rect 1548 987 1554 990
rect 156 950 162 953
rect 126 944 162 950
rect 810 950 816 953
rect 810 944 1584 950
rect 126 910 138 944
rect 1572 910 1584 944
rect 126 904 162 910
rect 156 901 162 904
rect 810 904 1584 910
rect 810 901 816 904
rect 894 864 900 867
rect 126 858 900 864
rect 1548 864 1554 867
rect 1548 858 1584 864
rect 126 824 138 858
rect 1572 824 1584 858
rect 126 818 900 824
rect 894 815 900 818
rect 1548 818 1584 824
rect 1548 815 1554 818
rect 156 778 162 781
rect 126 772 162 778
rect 810 778 816 781
rect 810 772 1584 778
rect 126 738 138 772
rect 1572 738 1584 772
rect 126 732 162 738
rect 156 729 162 732
rect 810 732 1584 738
rect 810 729 816 732
rect 894 692 900 695
rect 126 686 900 692
rect 1548 692 1554 695
rect 1548 686 1584 692
rect 126 652 138 686
rect 1572 652 1584 686
rect 126 646 900 652
rect 894 643 900 646
rect 1548 646 1584 652
rect 1548 643 1554 646
rect 156 606 162 609
rect 126 600 162 606
rect 810 606 816 609
rect 810 600 1584 606
rect 126 566 138 600
rect 1572 566 1584 600
rect 126 560 162 566
rect 156 557 162 560
rect 810 560 1584 566
rect 810 557 816 560
rect 894 520 900 523
rect 126 514 900 520
rect 1548 520 1554 523
rect 1548 514 1584 520
rect 126 480 138 514
rect 1572 480 1584 514
rect 126 474 900 480
rect 894 471 900 474
rect 1548 474 1584 480
rect 1548 471 1554 474
rect 156 434 162 437
rect 126 428 162 434
rect 810 434 816 437
rect 810 428 1584 434
rect 126 394 138 428
rect 1572 394 1584 428
rect 126 388 162 394
rect 156 385 162 388
rect 810 388 1584 394
rect 810 385 816 388
rect 894 348 900 351
rect 126 342 900 348
rect 1548 348 1554 351
rect 1548 342 1584 348
rect 126 308 138 342
rect 1572 308 1584 342
rect 126 302 900 308
rect 894 299 900 302
rect 1548 302 1584 308
rect 1548 299 1554 302
rect 156 262 162 265
rect 126 256 162 262
rect 810 262 816 265
rect 810 256 1584 262
rect 126 222 138 256
rect 1572 222 1584 256
rect 126 216 162 222
rect 156 213 162 216
rect 810 216 1584 222
rect 810 213 816 216
rect 894 176 900 179
rect 126 170 900 176
rect 1548 176 1554 179
rect 1548 170 1584 176
rect 126 136 138 170
rect 1572 136 1584 170
rect 1618 163 1672 169
rect 126 130 900 136
rect 894 127 900 130
rect 1548 130 1584 136
rect 1548 127 1554 130
rect 30 76 76 100
rect 1704 100 1710 100138
rect 1744 100 1750 100138
rect 1704 76 1750 100
rect 30 70 1750 76
rect 30 36 100 70
rect 1680 36 1750 70
rect 30 30 1750 36
<< via1 >>
rect 900 100102 1548 100111
rect 900 100068 1548 100102
rect 900 100059 1548 100068
rect 1618 100059 1672 100069
rect 162 100016 810 100025
rect 162 99982 810 100016
rect 162 99973 810 99982
rect 900 99930 1548 99939
rect 900 99896 1548 99930
rect 900 99887 1548 99896
rect 162 99844 810 99853
rect 162 99810 810 99844
rect 162 99801 810 99810
rect 900 99758 1548 99767
rect 900 99724 1548 99758
rect 900 99715 1548 99724
rect 162 99672 810 99681
rect 162 99638 810 99672
rect 162 99629 810 99638
rect 900 99586 1548 99595
rect 900 99552 1548 99586
rect 900 99543 1548 99552
rect 162 99500 810 99509
rect 162 99466 810 99500
rect 162 99457 810 99466
rect 900 99414 1548 99423
rect 900 99380 1548 99414
rect 900 99371 1548 99380
rect 162 99328 810 99337
rect 162 99294 810 99328
rect 162 99285 810 99294
rect 900 99242 1548 99251
rect 900 99208 1548 99242
rect 900 99199 1548 99208
rect 162 99156 810 99165
rect 162 99122 810 99156
rect 162 99113 810 99122
rect 900 99070 1548 99079
rect 900 99036 1548 99070
rect 900 99027 1548 99036
rect 162 98984 810 98993
rect 162 98950 810 98984
rect 162 98941 810 98950
rect 900 98898 1548 98907
rect 900 98864 1548 98898
rect 900 98855 1548 98864
rect 162 98812 810 98821
rect 162 98778 810 98812
rect 162 98769 810 98778
rect 900 98726 1548 98735
rect 900 98692 1548 98726
rect 900 98683 1548 98692
rect 162 98640 810 98649
rect 162 98606 810 98640
rect 162 98597 810 98606
rect 900 98554 1548 98563
rect 900 98520 1548 98554
rect 900 98511 1548 98520
rect 162 98468 810 98477
rect 162 98434 810 98468
rect 162 98425 810 98434
rect 900 98382 1548 98391
rect 900 98348 1548 98382
rect 900 98339 1548 98348
rect 162 98296 810 98305
rect 162 98262 810 98296
rect 162 98253 810 98262
rect 900 98210 1548 98219
rect 900 98176 1548 98210
rect 900 98167 1548 98176
rect 162 98124 810 98133
rect 162 98090 810 98124
rect 162 98081 810 98090
rect 900 98038 1548 98047
rect 900 98004 1548 98038
rect 900 97995 1548 98004
rect 162 97952 810 97961
rect 162 97918 810 97952
rect 162 97909 810 97918
rect 900 97866 1548 97875
rect 900 97832 1548 97866
rect 900 97823 1548 97832
rect 162 97780 810 97789
rect 162 97746 810 97780
rect 162 97737 810 97746
rect 900 97694 1548 97703
rect 900 97660 1548 97694
rect 900 97651 1548 97660
rect 162 97608 810 97617
rect 162 97574 810 97608
rect 162 97565 810 97574
rect 900 97522 1548 97531
rect 900 97488 1548 97522
rect 900 97479 1548 97488
rect 162 97436 810 97445
rect 162 97402 810 97436
rect 162 97393 810 97402
rect 900 97350 1548 97359
rect 900 97316 1548 97350
rect 900 97307 1548 97316
rect 162 97264 810 97273
rect 162 97230 810 97264
rect 162 97221 810 97230
rect 900 97178 1548 97187
rect 900 97144 1548 97178
rect 900 97135 1548 97144
rect 162 97092 810 97101
rect 162 97058 810 97092
rect 162 97049 810 97058
rect 900 97006 1548 97015
rect 900 96972 1548 97006
rect 900 96963 1548 96972
rect 162 96920 810 96929
rect 162 96886 810 96920
rect 162 96877 810 96886
rect 900 96834 1548 96843
rect 900 96800 1548 96834
rect 900 96791 1548 96800
rect 162 96748 810 96757
rect 162 96714 810 96748
rect 162 96705 810 96714
rect 900 96662 1548 96671
rect 900 96628 1548 96662
rect 900 96619 1548 96628
rect 162 96576 810 96585
rect 162 96542 810 96576
rect 162 96533 810 96542
rect 900 96490 1548 96499
rect 900 96456 1548 96490
rect 900 96447 1548 96456
rect 162 96404 810 96413
rect 162 96370 810 96404
rect 162 96361 810 96370
rect 900 96318 1548 96327
rect 900 96284 1548 96318
rect 900 96275 1548 96284
rect 162 96232 810 96241
rect 162 96198 810 96232
rect 162 96189 810 96198
rect 900 96146 1548 96155
rect 900 96112 1548 96146
rect 900 96103 1548 96112
rect 162 96060 810 96069
rect 162 96026 810 96060
rect 162 96017 810 96026
rect 900 95974 1548 95983
rect 900 95940 1548 95974
rect 900 95931 1548 95940
rect 162 95888 810 95897
rect 162 95854 810 95888
rect 162 95845 810 95854
rect 900 95802 1548 95811
rect 900 95768 1548 95802
rect 900 95759 1548 95768
rect 162 95716 810 95725
rect 162 95682 810 95716
rect 162 95673 810 95682
rect 900 95630 1548 95639
rect 900 95596 1548 95630
rect 900 95587 1548 95596
rect 162 95544 810 95553
rect 162 95510 810 95544
rect 162 95501 810 95510
rect 900 95458 1548 95467
rect 900 95424 1548 95458
rect 900 95415 1548 95424
rect 162 95372 810 95381
rect 162 95338 810 95372
rect 162 95329 810 95338
rect 900 95286 1548 95295
rect 900 95252 1548 95286
rect 900 95243 1548 95252
rect 162 95200 810 95209
rect 162 95166 810 95200
rect 162 95157 810 95166
rect 900 95114 1548 95123
rect 900 95080 1548 95114
rect 900 95071 1548 95080
rect 162 95028 810 95037
rect 162 94994 810 95028
rect 162 94985 810 94994
rect 900 94942 1548 94951
rect 900 94908 1548 94942
rect 900 94899 1548 94908
rect 162 94856 810 94865
rect 162 94822 810 94856
rect 162 94813 810 94822
rect 900 94770 1548 94779
rect 900 94736 1548 94770
rect 900 94727 1548 94736
rect 162 94684 810 94693
rect 162 94650 810 94684
rect 162 94641 810 94650
rect 900 94598 1548 94607
rect 900 94564 1548 94598
rect 900 94555 1548 94564
rect 162 94512 810 94521
rect 162 94478 810 94512
rect 162 94469 810 94478
rect 900 94426 1548 94435
rect 900 94392 1548 94426
rect 900 94383 1548 94392
rect 162 94340 810 94349
rect 162 94306 810 94340
rect 162 94297 810 94306
rect 900 94254 1548 94263
rect 900 94220 1548 94254
rect 900 94211 1548 94220
rect 162 94168 810 94177
rect 162 94134 810 94168
rect 162 94125 810 94134
rect 900 94082 1548 94091
rect 900 94048 1548 94082
rect 900 94039 1548 94048
rect 162 93996 810 94005
rect 162 93962 810 93996
rect 162 93953 810 93962
rect 900 93910 1548 93919
rect 900 93876 1548 93910
rect 900 93867 1548 93876
rect 162 93824 810 93833
rect 162 93790 810 93824
rect 162 93781 810 93790
rect 900 93738 1548 93747
rect 900 93704 1548 93738
rect 900 93695 1548 93704
rect 162 93652 810 93661
rect 162 93618 810 93652
rect 162 93609 810 93618
rect 900 93566 1548 93575
rect 900 93532 1548 93566
rect 900 93523 1548 93532
rect 162 93480 810 93489
rect 162 93446 810 93480
rect 162 93437 810 93446
rect 900 93394 1548 93403
rect 900 93360 1548 93394
rect 900 93351 1548 93360
rect 162 93308 810 93317
rect 162 93274 810 93308
rect 162 93265 810 93274
rect 900 93222 1548 93231
rect 900 93188 1548 93222
rect 900 93179 1548 93188
rect 162 93136 810 93145
rect 162 93102 810 93136
rect 162 93093 810 93102
rect 900 93050 1548 93059
rect 900 93016 1548 93050
rect 900 93007 1548 93016
rect 162 92964 810 92973
rect 162 92930 810 92964
rect 162 92921 810 92930
rect 900 92878 1548 92887
rect 900 92844 1548 92878
rect 900 92835 1548 92844
rect 162 92792 810 92801
rect 162 92758 810 92792
rect 162 92749 810 92758
rect 900 92706 1548 92715
rect 900 92672 1548 92706
rect 900 92663 1548 92672
rect 162 92620 810 92629
rect 162 92586 810 92620
rect 162 92577 810 92586
rect 900 92534 1548 92543
rect 900 92500 1548 92534
rect 900 92491 1548 92500
rect 162 92448 810 92457
rect 162 92414 810 92448
rect 162 92405 810 92414
rect 900 92362 1548 92371
rect 900 92328 1548 92362
rect 900 92319 1548 92328
rect 162 92276 810 92285
rect 162 92242 810 92276
rect 162 92233 810 92242
rect 900 92190 1548 92199
rect 900 92156 1548 92190
rect 900 92147 1548 92156
rect 162 92104 810 92113
rect 162 92070 810 92104
rect 162 92061 810 92070
rect 900 92018 1548 92027
rect 900 91984 1548 92018
rect 900 91975 1548 91984
rect 162 91932 810 91941
rect 162 91898 810 91932
rect 162 91889 810 91898
rect 900 91846 1548 91855
rect 900 91812 1548 91846
rect 900 91803 1548 91812
rect 162 91760 810 91769
rect 162 91726 810 91760
rect 162 91717 810 91726
rect 900 91674 1548 91683
rect 900 91640 1548 91674
rect 900 91631 1548 91640
rect 162 91588 810 91597
rect 162 91554 810 91588
rect 162 91545 810 91554
rect 900 91502 1548 91511
rect 900 91468 1548 91502
rect 900 91459 1548 91468
rect 162 91416 810 91425
rect 162 91382 810 91416
rect 162 91373 810 91382
rect 900 91330 1548 91339
rect 900 91296 1548 91330
rect 900 91287 1548 91296
rect 162 91244 810 91253
rect 162 91210 810 91244
rect 162 91201 810 91210
rect 900 91158 1548 91167
rect 900 91124 1548 91158
rect 900 91115 1548 91124
rect 162 91072 810 91081
rect 162 91038 810 91072
rect 162 91029 810 91038
rect 900 90986 1548 90995
rect 900 90952 1548 90986
rect 900 90943 1548 90952
rect 162 90900 810 90909
rect 162 90866 810 90900
rect 162 90857 810 90866
rect 900 90814 1548 90823
rect 900 90780 1548 90814
rect 900 90771 1548 90780
rect 162 90728 810 90737
rect 162 90694 810 90728
rect 162 90685 810 90694
rect 900 90642 1548 90651
rect 900 90608 1548 90642
rect 900 90599 1548 90608
rect 162 90556 810 90565
rect 162 90522 810 90556
rect 162 90513 810 90522
rect 900 90470 1548 90479
rect 900 90436 1548 90470
rect 900 90427 1548 90436
rect 162 90384 810 90393
rect 162 90350 810 90384
rect 162 90341 810 90350
rect 900 90298 1548 90307
rect 900 90264 1548 90298
rect 900 90255 1548 90264
rect 162 90212 810 90221
rect 162 90178 810 90212
rect 162 90169 810 90178
rect 900 90126 1548 90135
rect 900 90092 1548 90126
rect 900 90083 1548 90092
rect 162 90040 810 90049
rect 162 90006 810 90040
rect 162 89997 810 90006
rect 900 89954 1548 89963
rect 900 89920 1548 89954
rect 900 89911 1548 89920
rect 162 89868 810 89877
rect 162 89834 810 89868
rect 162 89825 810 89834
rect 900 89782 1548 89791
rect 900 89748 1548 89782
rect 900 89739 1548 89748
rect 162 89696 810 89705
rect 162 89662 810 89696
rect 162 89653 810 89662
rect 900 89610 1548 89619
rect 900 89576 1548 89610
rect 900 89567 1548 89576
rect 162 89524 810 89533
rect 162 89490 810 89524
rect 162 89481 810 89490
rect 900 89438 1548 89447
rect 900 89404 1548 89438
rect 900 89395 1548 89404
rect 162 89352 810 89361
rect 162 89318 810 89352
rect 162 89309 810 89318
rect 900 89266 1548 89275
rect 900 89232 1548 89266
rect 900 89223 1548 89232
rect 162 89180 810 89189
rect 162 89146 810 89180
rect 162 89137 810 89146
rect 900 89094 1548 89103
rect 900 89060 1548 89094
rect 900 89051 1548 89060
rect 162 89008 810 89017
rect 162 88974 810 89008
rect 162 88965 810 88974
rect 900 88922 1548 88931
rect 900 88888 1548 88922
rect 900 88879 1548 88888
rect 162 88836 810 88845
rect 162 88802 810 88836
rect 162 88793 810 88802
rect 900 88750 1548 88759
rect 900 88716 1548 88750
rect 900 88707 1548 88716
rect 162 88664 810 88673
rect 162 88630 810 88664
rect 162 88621 810 88630
rect 900 88578 1548 88587
rect 900 88544 1548 88578
rect 900 88535 1548 88544
rect 162 88492 810 88501
rect 162 88458 810 88492
rect 162 88449 810 88458
rect 900 88406 1548 88415
rect 900 88372 1548 88406
rect 900 88363 1548 88372
rect 162 88320 810 88329
rect 162 88286 810 88320
rect 162 88277 810 88286
rect 900 88234 1548 88243
rect 900 88200 1548 88234
rect 900 88191 1548 88200
rect 162 88148 810 88157
rect 162 88114 810 88148
rect 162 88105 810 88114
rect 900 88062 1548 88071
rect 900 88028 1548 88062
rect 900 88019 1548 88028
rect 162 87976 810 87985
rect 162 87942 810 87976
rect 162 87933 810 87942
rect 900 87890 1548 87899
rect 900 87856 1548 87890
rect 900 87847 1548 87856
rect 162 87804 810 87813
rect 162 87770 810 87804
rect 162 87761 810 87770
rect 900 87718 1548 87727
rect 900 87684 1548 87718
rect 900 87675 1548 87684
rect 162 87632 810 87641
rect 162 87598 810 87632
rect 162 87589 810 87598
rect 900 87546 1548 87555
rect 900 87512 1548 87546
rect 900 87503 1548 87512
rect 162 87460 810 87469
rect 162 87426 810 87460
rect 162 87417 810 87426
rect 900 87374 1548 87383
rect 900 87340 1548 87374
rect 900 87331 1548 87340
rect 162 87288 810 87297
rect 162 87254 810 87288
rect 162 87245 810 87254
rect 900 87202 1548 87211
rect 900 87168 1548 87202
rect 900 87159 1548 87168
rect 162 87116 810 87125
rect 162 87082 810 87116
rect 162 87073 810 87082
rect 900 87030 1548 87039
rect 900 86996 1548 87030
rect 900 86987 1548 86996
rect 162 86944 810 86953
rect 162 86910 810 86944
rect 162 86901 810 86910
rect 900 86858 1548 86867
rect 900 86824 1548 86858
rect 900 86815 1548 86824
rect 162 86772 810 86781
rect 162 86738 810 86772
rect 162 86729 810 86738
rect 900 86686 1548 86695
rect 900 86652 1548 86686
rect 900 86643 1548 86652
rect 162 86600 810 86609
rect 162 86566 810 86600
rect 162 86557 810 86566
rect 900 86514 1548 86523
rect 900 86480 1548 86514
rect 900 86471 1548 86480
rect 162 86428 810 86437
rect 162 86394 810 86428
rect 162 86385 810 86394
rect 900 86342 1548 86351
rect 900 86308 1548 86342
rect 900 86299 1548 86308
rect 162 86256 810 86265
rect 162 86222 810 86256
rect 162 86213 810 86222
rect 900 86170 1548 86179
rect 900 86136 1548 86170
rect 900 86127 1548 86136
rect 162 86084 810 86093
rect 162 86050 810 86084
rect 162 86041 810 86050
rect 900 85998 1548 86007
rect 900 85964 1548 85998
rect 900 85955 1548 85964
rect 162 85912 810 85921
rect 162 85878 810 85912
rect 162 85869 810 85878
rect 900 85826 1548 85835
rect 900 85792 1548 85826
rect 900 85783 1548 85792
rect 162 85740 810 85749
rect 162 85706 810 85740
rect 162 85697 810 85706
rect 900 85654 1548 85663
rect 900 85620 1548 85654
rect 900 85611 1548 85620
rect 162 85568 810 85577
rect 162 85534 810 85568
rect 162 85525 810 85534
rect 900 85482 1548 85491
rect 900 85448 1548 85482
rect 900 85439 1548 85448
rect 162 85396 810 85405
rect 162 85362 810 85396
rect 162 85353 810 85362
rect 900 85310 1548 85319
rect 900 85276 1548 85310
rect 900 85267 1548 85276
rect 162 85224 810 85233
rect 162 85190 810 85224
rect 162 85181 810 85190
rect 900 85138 1548 85147
rect 900 85104 1548 85138
rect 900 85095 1548 85104
rect 162 85052 810 85061
rect 162 85018 810 85052
rect 162 85009 810 85018
rect 900 84966 1548 84975
rect 900 84932 1548 84966
rect 900 84923 1548 84932
rect 162 84880 810 84889
rect 162 84846 810 84880
rect 162 84837 810 84846
rect 900 84794 1548 84803
rect 900 84760 1548 84794
rect 900 84751 1548 84760
rect 162 84708 810 84717
rect 162 84674 810 84708
rect 162 84665 810 84674
rect 900 84622 1548 84631
rect 900 84588 1548 84622
rect 900 84579 1548 84588
rect 162 84536 810 84545
rect 162 84502 810 84536
rect 162 84493 810 84502
rect 900 84450 1548 84459
rect 900 84416 1548 84450
rect 900 84407 1548 84416
rect 162 84364 810 84373
rect 162 84330 810 84364
rect 162 84321 810 84330
rect 900 84278 1548 84287
rect 900 84244 1548 84278
rect 900 84235 1548 84244
rect 162 84192 810 84201
rect 162 84158 810 84192
rect 162 84149 810 84158
rect 900 84106 1548 84115
rect 900 84072 1548 84106
rect 900 84063 1548 84072
rect 162 84020 810 84029
rect 162 83986 810 84020
rect 162 83977 810 83986
rect 900 83934 1548 83943
rect 900 83900 1548 83934
rect 900 83891 1548 83900
rect 162 83848 810 83857
rect 162 83814 810 83848
rect 162 83805 810 83814
rect 900 83762 1548 83771
rect 900 83728 1548 83762
rect 900 83719 1548 83728
rect 162 83676 810 83685
rect 162 83642 810 83676
rect 162 83633 810 83642
rect 900 83590 1548 83599
rect 900 83556 1548 83590
rect 900 83547 1548 83556
rect 162 83504 810 83513
rect 162 83470 810 83504
rect 162 83461 810 83470
rect 900 83418 1548 83427
rect 900 83384 1548 83418
rect 900 83375 1548 83384
rect 162 83332 810 83341
rect 162 83298 810 83332
rect 162 83289 810 83298
rect 900 83246 1548 83255
rect 900 83212 1548 83246
rect 900 83203 1548 83212
rect 162 83160 810 83169
rect 162 83126 810 83160
rect 162 83117 810 83126
rect 900 83074 1548 83083
rect 900 83040 1548 83074
rect 900 83031 1548 83040
rect 162 82988 810 82997
rect 162 82954 810 82988
rect 162 82945 810 82954
rect 900 82902 1548 82911
rect 900 82868 1548 82902
rect 900 82859 1548 82868
rect 162 82816 810 82825
rect 162 82782 810 82816
rect 162 82773 810 82782
rect 900 82730 1548 82739
rect 900 82696 1548 82730
rect 900 82687 1548 82696
rect 162 82644 810 82653
rect 162 82610 810 82644
rect 162 82601 810 82610
rect 900 82558 1548 82567
rect 900 82524 1548 82558
rect 900 82515 1548 82524
rect 162 82472 810 82481
rect 162 82438 810 82472
rect 162 82429 810 82438
rect 900 82386 1548 82395
rect 900 82352 1548 82386
rect 900 82343 1548 82352
rect 162 82300 810 82309
rect 162 82266 810 82300
rect 162 82257 810 82266
rect 900 82214 1548 82223
rect 900 82180 1548 82214
rect 900 82171 1548 82180
rect 162 82128 810 82137
rect 162 82094 810 82128
rect 162 82085 810 82094
rect 900 82042 1548 82051
rect 900 82008 1548 82042
rect 900 81999 1548 82008
rect 162 81956 810 81965
rect 162 81922 810 81956
rect 162 81913 810 81922
rect 900 81870 1548 81879
rect 900 81836 1548 81870
rect 900 81827 1548 81836
rect 162 81784 810 81793
rect 162 81750 810 81784
rect 162 81741 810 81750
rect 900 81698 1548 81707
rect 900 81664 1548 81698
rect 900 81655 1548 81664
rect 162 81612 810 81621
rect 162 81578 810 81612
rect 162 81569 810 81578
rect 900 81526 1548 81535
rect 900 81492 1548 81526
rect 900 81483 1548 81492
rect 162 81440 810 81449
rect 162 81406 810 81440
rect 162 81397 810 81406
rect 900 81354 1548 81363
rect 900 81320 1548 81354
rect 900 81311 1548 81320
rect 162 81268 810 81277
rect 162 81234 810 81268
rect 162 81225 810 81234
rect 900 81182 1548 81191
rect 900 81148 1548 81182
rect 900 81139 1548 81148
rect 162 81096 810 81105
rect 162 81062 810 81096
rect 162 81053 810 81062
rect 900 81010 1548 81019
rect 900 80976 1548 81010
rect 900 80967 1548 80976
rect 162 80924 810 80933
rect 162 80890 810 80924
rect 162 80881 810 80890
rect 900 80838 1548 80847
rect 900 80804 1548 80838
rect 900 80795 1548 80804
rect 162 80752 810 80761
rect 162 80718 810 80752
rect 162 80709 810 80718
rect 900 80666 1548 80675
rect 900 80632 1548 80666
rect 900 80623 1548 80632
rect 162 80580 810 80589
rect 162 80546 810 80580
rect 162 80537 810 80546
rect 900 80494 1548 80503
rect 900 80460 1548 80494
rect 900 80451 1548 80460
rect 162 80408 810 80417
rect 162 80374 810 80408
rect 162 80365 810 80374
rect 900 80322 1548 80331
rect 900 80288 1548 80322
rect 900 80279 1548 80288
rect 162 80236 810 80245
rect 162 80202 810 80236
rect 162 80193 810 80202
rect 900 80150 1548 80159
rect 900 80116 1548 80150
rect 900 80107 1548 80116
rect 162 80064 810 80073
rect 162 80030 810 80064
rect 162 80021 810 80030
rect 900 79978 1548 79987
rect 900 79944 1548 79978
rect 900 79935 1548 79944
rect 162 79892 810 79901
rect 162 79858 810 79892
rect 162 79849 810 79858
rect 900 79806 1548 79815
rect 900 79772 1548 79806
rect 900 79763 1548 79772
rect 162 79720 810 79729
rect 162 79686 810 79720
rect 162 79677 810 79686
rect 900 79634 1548 79643
rect 900 79600 1548 79634
rect 900 79591 1548 79600
rect 162 79548 810 79557
rect 162 79514 810 79548
rect 162 79505 810 79514
rect 900 79462 1548 79471
rect 900 79428 1548 79462
rect 900 79419 1548 79428
rect 162 79376 810 79385
rect 162 79342 810 79376
rect 162 79333 810 79342
rect 900 79290 1548 79299
rect 900 79256 1548 79290
rect 900 79247 1548 79256
rect 162 79204 810 79213
rect 162 79170 810 79204
rect 162 79161 810 79170
rect 900 79118 1548 79127
rect 900 79084 1548 79118
rect 900 79075 1548 79084
rect 162 79032 810 79041
rect 162 78998 810 79032
rect 162 78989 810 78998
rect 900 78946 1548 78955
rect 900 78912 1548 78946
rect 900 78903 1548 78912
rect 162 78860 810 78869
rect 162 78826 810 78860
rect 162 78817 810 78826
rect 900 78774 1548 78783
rect 900 78740 1548 78774
rect 900 78731 1548 78740
rect 162 78688 810 78697
rect 162 78654 810 78688
rect 162 78645 810 78654
rect 900 78602 1548 78611
rect 900 78568 1548 78602
rect 900 78559 1548 78568
rect 162 78516 810 78525
rect 162 78482 810 78516
rect 162 78473 810 78482
rect 900 78430 1548 78439
rect 900 78396 1548 78430
rect 900 78387 1548 78396
rect 162 78344 810 78353
rect 162 78310 810 78344
rect 162 78301 810 78310
rect 900 78258 1548 78267
rect 900 78224 1548 78258
rect 900 78215 1548 78224
rect 162 78172 810 78181
rect 162 78138 810 78172
rect 162 78129 810 78138
rect 900 78086 1548 78095
rect 900 78052 1548 78086
rect 900 78043 1548 78052
rect 162 78000 810 78009
rect 162 77966 810 78000
rect 162 77957 810 77966
rect 900 77914 1548 77923
rect 900 77880 1548 77914
rect 900 77871 1548 77880
rect 162 77828 810 77837
rect 162 77794 810 77828
rect 162 77785 810 77794
rect 900 77742 1548 77751
rect 900 77708 1548 77742
rect 900 77699 1548 77708
rect 162 77656 810 77665
rect 162 77622 810 77656
rect 162 77613 810 77622
rect 900 77570 1548 77579
rect 900 77536 1548 77570
rect 900 77527 1548 77536
rect 162 77484 810 77493
rect 162 77450 810 77484
rect 162 77441 810 77450
rect 900 77398 1548 77407
rect 900 77364 1548 77398
rect 900 77355 1548 77364
rect 162 77312 810 77321
rect 162 77278 810 77312
rect 162 77269 810 77278
rect 900 77226 1548 77235
rect 900 77192 1548 77226
rect 900 77183 1548 77192
rect 162 77140 810 77149
rect 162 77106 810 77140
rect 162 77097 810 77106
rect 900 77054 1548 77063
rect 900 77020 1548 77054
rect 900 77011 1548 77020
rect 162 76968 810 76977
rect 162 76934 810 76968
rect 162 76925 810 76934
rect 900 76882 1548 76891
rect 900 76848 1548 76882
rect 900 76839 1548 76848
rect 162 76796 810 76805
rect 162 76762 810 76796
rect 162 76753 810 76762
rect 900 76710 1548 76719
rect 900 76676 1548 76710
rect 900 76667 1548 76676
rect 162 76624 810 76633
rect 162 76590 810 76624
rect 162 76581 810 76590
rect 900 76538 1548 76547
rect 900 76504 1548 76538
rect 900 76495 1548 76504
rect 162 76452 810 76461
rect 162 76418 810 76452
rect 162 76409 810 76418
rect 900 76366 1548 76375
rect 900 76332 1548 76366
rect 900 76323 1548 76332
rect 162 76280 810 76289
rect 162 76246 810 76280
rect 162 76237 810 76246
rect 900 76194 1548 76203
rect 900 76160 1548 76194
rect 900 76151 1548 76160
rect 162 76108 810 76117
rect 162 76074 810 76108
rect 162 76065 810 76074
rect 900 76022 1548 76031
rect 900 75988 1548 76022
rect 900 75979 1548 75988
rect 162 75936 810 75945
rect 162 75902 810 75936
rect 162 75893 810 75902
rect 900 75850 1548 75859
rect 900 75816 1548 75850
rect 900 75807 1548 75816
rect 162 75764 810 75773
rect 162 75730 810 75764
rect 162 75721 810 75730
rect 900 75678 1548 75687
rect 900 75644 1548 75678
rect 900 75635 1548 75644
rect 162 75592 810 75601
rect 162 75558 810 75592
rect 162 75549 810 75558
rect 900 75506 1548 75515
rect 900 75472 1548 75506
rect 900 75463 1548 75472
rect 162 75420 810 75429
rect 162 75386 810 75420
rect 162 75377 810 75386
rect 900 75334 1548 75343
rect 900 75300 1548 75334
rect 900 75291 1548 75300
rect 162 75248 810 75257
rect 162 75214 810 75248
rect 162 75205 810 75214
rect 900 75162 1548 75171
rect 900 75128 1548 75162
rect 900 75119 1548 75128
rect 162 75076 810 75085
rect 162 75042 810 75076
rect 162 75033 810 75042
rect 900 74990 1548 74999
rect 900 74956 1548 74990
rect 900 74947 1548 74956
rect 162 74904 810 74913
rect 162 74870 810 74904
rect 162 74861 810 74870
rect 900 74818 1548 74827
rect 900 74784 1548 74818
rect 900 74775 1548 74784
rect 162 74732 810 74741
rect 162 74698 810 74732
rect 162 74689 810 74698
rect 900 74646 1548 74655
rect 900 74612 1548 74646
rect 900 74603 1548 74612
rect 162 74560 810 74569
rect 162 74526 810 74560
rect 162 74517 810 74526
rect 900 74474 1548 74483
rect 900 74440 1548 74474
rect 900 74431 1548 74440
rect 162 74388 810 74397
rect 162 74354 810 74388
rect 162 74345 810 74354
rect 900 74302 1548 74311
rect 900 74268 1548 74302
rect 900 74259 1548 74268
rect 162 74216 810 74225
rect 162 74182 810 74216
rect 162 74173 810 74182
rect 900 74130 1548 74139
rect 900 74096 1548 74130
rect 900 74087 1548 74096
rect 162 74044 810 74053
rect 162 74010 810 74044
rect 162 74001 810 74010
rect 900 73958 1548 73967
rect 900 73924 1548 73958
rect 900 73915 1548 73924
rect 162 73872 810 73881
rect 162 73838 810 73872
rect 162 73829 810 73838
rect 900 73786 1548 73795
rect 900 73752 1548 73786
rect 900 73743 1548 73752
rect 162 73700 810 73709
rect 162 73666 810 73700
rect 162 73657 810 73666
rect 900 73614 1548 73623
rect 900 73580 1548 73614
rect 900 73571 1548 73580
rect 162 73528 810 73537
rect 162 73494 810 73528
rect 162 73485 810 73494
rect 900 73442 1548 73451
rect 900 73408 1548 73442
rect 900 73399 1548 73408
rect 162 73356 810 73365
rect 162 73322 810 73356
rect 162 73313 810 73322
rect 900 73270 1548 73279
rect 900 73236 1548 73270
rect 900 73227 1548 73236
rect 162 73184 810 73193
rect 162 73150 810 73184
rect 162 73141 810 73150
rect 900 73098 1548 73107
rect 900 73064 1548 73098
rect 900 73055 1548 73064
rect 162 73012 810 73021
rect 162 72978 810 73012
rect 162 72969 810 72978
rect 900 72926 1548 72935
rect 900 72892 1548 72926
rect 900 72883 1548 72892
rect 162 72840 810 72849
rect 162 72806 810 72840
rect 162 72797 810 72806
rect 900 72754 1548 72763
rect 900 72720 1548 72754
rect 900 72711 1548 72720
rect 162 72668 810 72677
rect 162 72634 810 72668
rect 162 72625 810 72634
rect 900 72582 1548 72591
rect 900 72548 1548 72582
rect 900 72539 1548 72548
rect 162 72496 810 72505
rect 162 72462 810 72496
rect 162 72453 810 72462
rect 900 72410 1548 72419
rect 900 72376 1548 72410
rect 900 72367 1548 72376
rect 162 72324 810 72333
rect 162 72290 810 72324
rect 162 72281 810 72290
rect 900 72238 1548 72247
rect 900 72204 1548 72238
rect 900 72195 1548 72204
rect 162 72152 810 72161
rect 162 72118 810 72152
rect 162 72109 810 72118
rect 900 72066 1548 72075
rect 900 72032 1548 72066
rect 900 72023 1548 72032
rect 162 71980 810 71989
rect 162 71946 810 71980
rect 162 71937 810 71946
rect 900 71894 1548 71903
rect 900 71860 1548 71894
rect 900 71851 1548 71860
rect 162 71808 810 71817
rect 162 71774 810 71808
rect 162 71765 810 71774
rect 900 71722 1548 71731
rect 900 71688 1548 71722
rect 900 71679 1548 71688
rect 162 71636 810 71645
rect 162 71602 810 71636
rect 162 71593 810 71602
rect 900 71550 1548 71559
rect 900 71516 1548 71550
rect 900 71507 1548 71516
rect 162 71464 810 71473
rect 162 71430 810 71464
rect 162 71421 810 71430
rect 900 71378 1548 71387
rect 900 71344 1548 71378
rect 900 71335 1548 71344
rect 162 71292 810 71301
rect 162 71258 810 71292
rect 162 71249 810 71258
rect 900 71206 1548 71215
rect 900 71172 1548 71206
rect 900 71163 1548 71172
rect 162 71120 810 71129
rect 162 71086 810 71120
rect 162 71077 810 71086
rect 900 71034 1548 71043
rect 900 71000 1548 71034
rect 900 70991 1548 71000
rect 162 70948 810 70957
rect 162 70914 810 70948
rect 162 70905 810 70914
rect 900 70862 1548 70871
rect 900 70828 1548 70862
rect 900 70819 1548 70828
rect 162 70776 810 70785
rect 162 70742 810 70776
rect 162 70733 810 70742
rect 900 70690 1548 70699
rect 900 70656 1548 70690
rect 900 70647 1548 70656
rect 162 70604 810 70613
rect 162 70570 810 70604
rect 162 70561 810 70570
rect 900 70518 1548 70527
rect 900 70484 1548 70518
rect 900 70475 1548 70484
rect 162 70432 810 70441
rect 162 70398 810 70432
rect 162 70389 810 70398
rect 900 70346 1548 70355
rect 900 70312 1548 70346
rect 900 70303 1548 70312
rect 162 70260 810 70269
rect 162 70226 810 70260
rect 162 70217 810 70226
rect 900 70174 1548 70183
rect 900 70140 1548 70174
rect 900 70131 1548 70140
rect 162 70088 810 70097
rect 162 70054 810 70088
rect 162 70045 810 70054
rect 900 70002 1548 70011
rect 900 69968 1548 70002
rect 900 69959 1548 69968
rect 162 69916 810 69925
rect 162 69882 810 69916
rect 162 69873 810 69882
rect 900 69830 1548 69839
rect 900 69796 1548 69830
rect 900 69787 1548 69796
rect 162 69744 810 69753
rect 162 69710 810 69744
rect 162 69701 810 69710
rect 900 69658 1548 69667
rect 900 69624 1548 69658
rect 900 69615 1548 69624
rect 162 69572 810 69581
rect 162 69538 810 69572
rect 162 69529 810 69538
rect 900 69486 1548 69495
rect 900 69452 1548 69486
rect 900 69443 1548 69452
rect 162 69400 810 69409
rect 162 69366 810 69400
rect 162 69357 810 69366
rect 900 69314 1548 69323
rect 900 69280 1548 69314
rect 900 69271 1548 69280
rect 162 69228 810 69237
rect 162 69194 810 69228
rect 162 69185 810 69194
rect 900 69142 1548 69151
rect 900 69108 1548 69142
rect 900 69099 1548 69108
rect 162 69056 810 69065
rect 162 69022 810 69056
rect 162 69013 810 69022
rect 900 68970 1548 68979
rect 900 68936 1548 68970
rect 900 68927 1548 68936
rect 162 68884 810 68893
rect 162 68850 810 68884
rect 162 68841 810 68850
rect 900 68798 1548 68807
rect 900 68764 1548 68798
rect 900 68755 1548 68764
rect 162 68712 810 68721
rect 162 68678 810 68712
rect 162 68669 810 68678
rect 900 68626 1548 68635
rect 900 68592 1548 68626
rect 900 68583 1548 68592
rect 162 68540 810 68549
rect 162 68506 810 68540
rect 162 68497 810 68506
rect 900 68454 1548 68463
rect 900 68420 1548 68454
rect 900 68411 1548 68420
rect 162 68368 810 68377
rect 162 68334 810 68368
rect 162 68325 810 68334
rect 900 68282 1548 68291
rect 900 68248 1548 68282
rect 900 68239 1548 68248
rect 162 68196 810 68205
rect 162 68162 810 68196
rect 162 68153 810 68162
rect 900 68110 1548 68119
rect 900 68076 1548 68110
rect 900 68067 1548 68076
rect 162 68024 810 68033
rect 162 67990 810 68024
rect 162 67981 810 67990
rect 900 67938 1548 67947
rect 900 67904 1548 67938
rect 900 67895 1548 67904
rect 162 67852 810 67861
rect 162 67818 810 67852
rect 162 67809 810 67818
rect 900 67766 1548 67775
rect 900 67732 1548 67766
rect 900 67723 1548 67732
rect 162 67680 810 67689
rect 162 67646 810 67680
rect 162 67637 810 67646
rect 900 67594 1548 67603
rect 900 67560 1548 67594
rect 900 67551 1548 67560
rect 162 67508 810 67517
rect 162 67474 810 67508
rect 162 67465 810 67474
rect 900 67422 1548 67431
rect 900 67388 1548 67422
rect 900 67379 1548 67388
rect 162 67336 810 67345
rect 162 67302 810 67336
rect 162 67293 810 67302
rect 900 67250 1548 67259
rect 900 67216 1548 67250
rect 900 67207 1548 67216
rect 162 67164 810 67173
rect 162 67130 810 67164
rect 162 67121 810 67130
rect 900 67078 1548 67087
rect 900 67044 1548 67078
rect 900 67035 1548 67044
rect 162 66992 810 67001
rect 162 66958 810 66992
rect 162 66949 810 66958
rect 900 66906 1548 66915
rect 900 66872 1548 66906
rect 900 66863 1548 66872
rect 162 66820 810 66829
rect 162 66786 810 66820
rect 162 66777 810 66786
rect 900 66734 1548 66743
rect 900 66700 1548 66734
rect 900 66691 1548 66700
rect 162 66648 810 66657
rect 162 66614 810 66648
rect 162 66605 810 66614
rect 900 66562 1548 66571
rect 900 66528 1548 66562
rect 900 66519 1548 66528
rect 162 66476 810 66485
rect 162 66442 810 66476
rect 162 66433 810 66442
rect 900 66390 1548 66399
rect 900 66356 1548 66390
rect 900 66347 1548 66356
rect 162 66304 810 66313
rect 162 66270 810 66304
rect 162 66261 810 66270
rect 900 66218 1548 66227
rect 900 66184 1548 66218
rect 900 66175 1548 66184
rect 162 66132 810 66141
rect 162 66098 810 66132
rect 162 66089 810 66098
rect 900 66046 1548 66055
rect 900 66012 1548 66046
rect 900 66003 1548 66012
rect 162 65960 810 65969
rect 162 65926 810 65960
rect 162 65917 810 65926
rect 900 65874 1548 65883
rect 900 65840 1548 65874
rect 900 65831 1548 65840
rect 162 65788 810 65797
rect 162 65754 810 65788
rect 162 65745 810 65754
rect 900 65702 1548 65711
rect 900 65668 1548 65702
rect 900 65659 1548 65668
rect 162 65616 810 65625
rect 162 65582 810 65616
rect 162 65573 810 65582
rect 900 65530 1548 65539
rect 900 65496 1548 65530
rect 900 65487 1548 65496
rect 162 65444 810 65453
rect 162 65410 810 65444
rect 162 65401 810 65410
rect 900 65358 1548 65367
rect 900 65324 1548 65358
rect 900 65315 1548 65324
rect 162 65272 810 65281
rect 162 65238 810 65272
rect 162 65229 810 65238
rect 900 65186 1548 65195
rect 900 65152 1548 65186
rect 900 65143 1548 65152
rect 162 65100 810 65109
rect 162 65066 810 65100
rect 162 65057 810 65066
rect 900 65014 1548 65023
rect 900 64980 1548 65014
rect 900 64971 1548 64980
rect 162 64928 810 64937
rect 162 64894 810 64928
rect 162 64885 810 64894
rect 900 64842 1548 64851
rect 900 64808 1548 64842
rect 900 64799 1548 64808
rect 162 64756 810 64765
rect 162 64722 810 64756
rect 162 64713 810 64722
rect 900 64670 1548 64679
rect 900 64636 1548 64670
rect 900 64627 1548 64636
rect 162 64584 810 64593
rect 162 64550 810 64584
rect 162 64541 810 64550
rect 900 64498 1548 64507
rect 900 64464 1548 64498
rect 900 64455 1548 64464
rect 162 64412 810 64421
rect 162 64378 810 64412
rect 162 64369 810 64378
rect 900 64326 1548 64335
rect 900 64292 1548 64326
rect 900 64283 1548 64292
rect 162 64240 810 64249
rect 162 64206 810 64240
rect 162 64197 810 64206
rect 900 64154 1548 64163
rect 900 64120 1548 64154
rect 900 64111 1548 64120
rect 162 64068 810 64077
rect 162 64034 810 64068
rect 162 64025 810 64034
rect 900 63982 1548 63991
rect 900 63948 1548 63982
rect 900 63939 1548 63948
rect 162 63896 810 63905
rect 162 63862 810 63896
rect 162 63853 810 63862
rect 900 63810 1548 63819
rect 900 63776 1548 63810
rect 900 63767 1548 63776
rect 162 63724 810 63733
rect 162 63690 810 63724
rect 162 63681 810 63690
rect 900 63638 1548 63647
rect 900 63604 1548 63638
rect 900 63595 1548 63604
rect 162 63552 810 63561
rect 162 63518 810 63552
rect 162 63509 810 63518
rect 900 63466 1548 63475
rect 900 63432 1548 63466
rect 900 63423 1548 63432
rect 162 63380 810 63389
rect 162 63346 810 63380
rect 162 63337 810 63346
rect 900 63294 1548 63303
rect 900 63260 1548 63294
rect 900 63251 1548 63260
rect 162 63208 810 63217
rect 162 63174 810 63208
rect 162 63165 810 63174
rect 900 63122 1548 63131
rect 900 63088 1548 63122
rect 900 63079 1548 63088
rect 162 63036 810 63045
rect 162 63002 810 63036
rect 162 62993 810 63002
rect 900 62950 1548 62959
rect 900 62916 1548 62950
rect 900 62907 1548 62916
rect 162 62864 810 62873
rect 162 62830 810 62864
rect 162 62821 810 62830
rect 900 62778 1548 62787
rect 900 62744 1548 62778
rect 900 62735 1548 62744
rect 162 62692 810 62701
rect 162 62658 810 62692
rect 162 62649 810 62658
rect 900 62606 1548 62615
rect 900 62572 1548 62606
rect 900 62563 1548 62572
rect 162 62520 810 62529
rect 162 62486 810 62520
rect 162 62477 810 62486
rect 900 62434 1548 62443
rect 900 62400 1548 62434
rect 900 62391 1548 62400
rect 162 62348 810 62357
rect 162 62314 810 62348
rect 162 62305 810 62314
rect 900 62262 1548 62271
rect 900 62228 1548 62262
rect 900 62219 1548 62228
rect 162 62176 810 62185
rect 162 62142 810 62176
rect 162 62133 810 62142
rect 900 62090 1548 62099
rect 900 62056 1548 62090
rect 900 62047 1548 62056
rect 162 62004 810 62013
rect 162 61970 810 62004
rect 162 61961 810 61970
rect 900 61918 1548 61927
rect 900 61884 1548 61918
rect 900 61875 1548 61884
rect 162 61832 810 61841
rect 162 61798 810 61832
rect 162 61789 810 61798
rect 900 61746 1548 61755
rect 900 61712 1548 61746
rect 900 61703 1548 61712
rect 162 61660 810 61669
rect 162 61626 810 61660
rect 162 61617 810 61626
rect 900 61574 1548 61583
rect 900 61540 1548 61574
rect 900 61531 1548 61540
rect 162 61488 810 61497
rect 162 61454 810 61488
rect 162 61445 810 61454
rect 900 61402 1548 61411
rect 900 61368 1548 61402
rect 900 61359 1548 61368
rect 162 61316 810 61325
rect 162 61282 810 61316
rect 162 61273 810 61282
rect 900 61230 1548 61239
rect 900 61196 1548 61230
rect 900 61187 1548 61196
rect 162 61144 810 61153
rect 162 61110 810 61144
rect 162 61101 810 61110
rect 900 61058 1548 61067
rect 900 61024 1548 61058
rect 900 61015 1548 61024
rect 162 60972 810 60981
rect 162 60938 810 60972
rect 162 60929 810 60938
rect 900 60886 1548 60895
rect 900 60852 1548 60886
rect 900 60843 1548 60852
rect 162 60800 810 60809
rect 162 60766 810 60800
rect 162 60757 810 60766
rect 900 60714 1548 60723
rect 900 60680 1548 60714
rect 900 60671 1548 60680
rect 162 60628 810 60637
rect 162 60594 810 60628
rect 162 60585 810 60594
rect 900 60542 1548 60551
rect 900 60508 1548 60542
rect 900 60499 1548 60508
rect 162 60456 810 60465
rect 162 60422 810 60456
rect 162 60413 810 60422
rect 900 60370 1548 60379
rect 900 60336 1548 60370
rect 900 60327 1548 60336
rect 162 60284 810 60293
rect 162 60250 810 60284
rect 162 60241 810 60250
rect 900 60198 1548 60207
rect 900 60164 1548 60198
rect 900 60155 1548 60164
rect 162 60112 810 60121
rect 162 60078 810 60112
rect 162 60069 810 60078
rect 900 60026 1548 60035
rect 900 59992 1548 60026
rect 900 59983 1548 59992
rect 162 59940 810 59949
rect 162 59906 810 59940
rect 162 59897 810 59906
rect 900 59854 1548 59863
rect 900 59820 1548 59854
rect 900 59811 1548 59820
rect 162 59768 810 59777
rect 162 59734 810 59768
rect 162 59725 810 59734
rect 900 59682 1548 59691
rect 900 59648 1548 59682
rect 900 59639 1548 59648
rect 162 59596 810 59605
rect 162 59562 810 59596
rect 162 59553 810 59562
rect 900 59510 1548 59519
rect 900 59476 1548 59510
rect 900 59467 1548 59476
rect 162 59424 810 59433
rect 162 59390 810 59424
rect 162 59381 810 59390
rect 900 59338 1548 59347
rect 900 59304 1548 59338
rect 900 59295 1548 59304
rect 162 59252 810 59261
rect 162 59218 810 59252
rect 162 59209 810 59218
rect 900 59166 1548 59175
rect 900 59132 1548 59166
rect 900 59123 1548 59132
rect 162 59080 810 59089
rect 162 59046 810 59080
rect 162 59037 810 59046
rect 900 58994 1548 59003
rect 900 58960 1548 58994
rect 900 58951 1548 58960
rect 162 58908 810 58917
rect 162 58874 810 58908
rect 162 58865 810 58874
rect 900 58822 1548 58831
rect 900 58788 1548 58822
rect 900 58779 1548 58788
rect 162 58736 810 58745
rect 162 58702 810 58736
rect 162 58693 810 58702
rect 900 58650 1548 58659
rect 900 58616 1548 58650
rect 900 58607 1548 58616
rect 162 58564 810 58573
rect 162 58530 810 58564
rect 162 58521 810 58530
rect 900 58478 1548 58487
rect 900 58444 1548 58478
rect 900 58435 1548 58444
rect 162 58392 810 58401
rect 162 58358 810 58392
rect 162 58349 810 58358
rect 900 58306 1548 58315
rect 900 58272 1548 58306
rect 900 58263 1548 58272
rect 162 58220 810 58229
rect 162 58186 810 58220
rect 162 58177 810 58186
rect 900 58134 1548 58143
rect 900 58100 1548 58134
rect 900 58091 1548 58100
rect 162 58048 810 58057
rect 162 58014 810 58048
rect 162 58005 810 58014
rect 900 57962 1548 57971
rect 900 57928 1548 57962
rect 900 57919 1548 57928
rect 162 57876 810 57885
rect 162 57842 810 57876
rect 162 57833 810 57842
rect 900 57790 1548 57799
rect 900 57756 1548 57790
rect 900 57747 1548 57756
rect 162 57704 810 57713
rect 162 57670 810 57704
rect 162 57661 810 57670
rect 900 57618 1548 57627
rect 900 57584 1548 57618
rect 900 57575 1548 57584
rect 162 57532 810 57541
rect 162 57498 810 57532
rect 162 57489 810 57498
rect 900 57446 1548 57455
rect 900 57412 1548 57446
rect 900 57403 1548 57412
rect 162 57360 810 57369
rect 162 57326 810 57360
rect 162 57317 810 57326
rect 900 57274 1548 57283
rect 900 57240 1548 57274
rect 900 57231 1548 57240
rect 162 57188 810 57197
rect 162 57154 810 57188
rect 162 57145 810 57154
rect 900 57102 1548 57111
rect 900 57068 1548 57102
rect 900 57059 1548 57068
rect 162 57016 810 57025
rect 162 56982 810 57016
rect 162 56973 810 56982
rect 900 56930 1548 56939
rect 900 56896 1548 56930
rect 900 56887 1548 56896
rect 162 56844 810 56853
rect 162 56810 810 56844
rect 162 56801 810 56810
rect 900 56758 1548 56767
rect 900 56724 1548 56758
rect 900 56715 1548 56724
rect 162 56672 810 56681
rect 162 56638 810 56672
rect 162 56629 810 56638
rect 900 56586 1548 56595
rect 900 56552 1548 56586
rect 900 56543 1548 56552
rect 162 56500 810 56509
rect 162 56466 810 56500
rect 162 56457 810 56466
rect 900 56414 1548 56423
rect 900 56380 1548 56414
rect 900 56371 1548 56380
rect 162 56328 810 56337
rect 162 56294 810 56328
rect 162 56285 810 56294
rect 900 56242 1548 56251
rect 900 56208 1548 56242
rect 900 56199 1548 56208
rect 162 56156 810 56165
rect 162 56122 810 56156
rect 162 56113 810 56122
rect 900 56070 1548 56079
rect 900 56036 1548 56070
rect 900 56027 1548 56036
rect 162 55984 810 55993
rect 162 55950 810 55984
rect 162 55941 810 55950
rect 900 55898 1548 55907
rect 900 55864 1548 55898
rect 900 55855 1548 55864
rect 162 55812 810 55821
rect 162 55778 810 55812
rect 162 55769 810 55778
rect 900 55726 1548 55735
rect 900 55692 1548 55726
rect 900 55683 1548 55692
rect 162 55640 810 55649
rect 162 55606 810 55640
rect 162 55597 810 55606
rect 900 55554 1548 55563
rect 900 55520 1548 55554
rect 900 55511 1548 55520
rect 162 55468 810 55477
rect 162 55434 810 55468
rect 162 55425 810 55434
rect 900 55382 1548 55391
rect 900 55348 1548 55382
rect 900 55339 1548 55348
rect 162 55296 810 55305
rect 162 55262 810 55296
rect 162 55253 810 55262
rect 900 55210 1548 55219
rect 900 55176 1548 55210
rect 900 55167 1548 55176
rect 162 55124 810 55133
rect 162 55090 810 55124
rect 162 55081 810 55090
rect 900 55038 1548 55047
rect 900 55004 1548 55038
rect 900 54995 1548 55004
rect 162 54952 810 54961
rect 162 54918 810 54952
rect 162 54909 810 54918
rect 900 54866 1548 54875
rect 900 54832 1548 54866
rect 900 54823 1548 54832
rect 162 54780 810 54789
rect 162 54746 810 54780
rect 162 54737 810 54746
rect 900 54694 1548 54703
rect 900 54660 1548 54694
rect 900 54651 1548 54660
rect 162 54608 810 54617
rect 162 54574 810 54608
rect 162 54565 810 54574
rect 900 54522 1548 54531
rect 900 54488 1548 54522
rect 900 54479 1548 54488
rect 162 54436 810 54445
rect 162 54402 810 54436
rect 162 54393 810 54402
rect 900 54350 1548 54359
rect 900 54316 1548 54350
rect 900 54307 1548 54316
rect 162 54264 810 54273
rect 162 54230 810 54264
rect 162 54221 810 54230
rect 900 54178 1548 54187
rect 900 54144 1548 54178
rect 900 54135 1548 54144
rect 162 54092 810 54101
rect 162 54058 810 54092
rect 162 54049 810 54058
rect 900 54006 1548 54015
rect 900 53972 1548 54006
rect 900 53963 1548 53972
rect 162 53920 810 53929
rect 162 53886 810 53920
rect 162 53877 810 53886
rect 900 53834 1548 53843
rect 900 53800 1548 53834
rect 900 53791 1548 53800
rect 162 53748 810 53757
rect 162 53714 810 53748
rect 162 53705 810 53714
rect 900 53662 1548 53671
rect 900 53628 1548 53662
rect 900 53619 1548 53628
rect 162 53576 810 53585
rect 162 53542 810 53576
rect 162 53533 810 53542
rect 900 53490 1548 53499
rect 900 53456 1548 53490
rect 900 53447 1548 53456
rect 162 53404 810 53413
rect 162 53370 810 53404
rect 162 53361 810 53370
rect 900 53318 1548 53327
rect 900 53284 1548 53318
rect 900 53275 1548 53284
rect 162 53232 810 53241
rect 162 53198 810 53232
rect 162 53189 810 53198
rect 900 53146 1548 53155
rect 900 53112 1548 53146
rect 900 53103 1548 53112
rect 162 53060 810 53069
rect 162 53026 810 53060
rect 162 53017 810 53026
rect 900 52974 1548 52983
rect 900 52940 1548 52974
rect 900 52931 1548 52940
rect 162 52888 810 52897
rect 162 52854 810 52888
rect 162 52845 810 52854
rect 900 52802 1548 52811
rect 900 52768 1548 52802
rect 900 52759 1548 52768
rect 162 52716 810 52725
rect 162 52682 810 52716
rect 162 52673 810 52682
rect 900 52630 1548 52639
rect 900 52596 1548 52630
rect 900 52587 1548 52596
rect 162 52544 810 52553
rect 162 52510 810 52544
rect 162 52501 810 52510
rect 900 52458 1548 52467
rect 900 52424 1548 52458
rect 900 52415 1548 52424
rect 162 52372 810 52381
rect 162 52338 810 52372
rect 162 52329 810 52338
rect 900 52286 1548 52295
rect 900 52252 1548 52286
rect 900 52243 1548 52252
rect 162 52200 810 52209
rect 162 52166 810 52200
rect 162 52157 810 52166
rect 900 52114 1548 52123
rect 900 52080 1548 52114
rect 900 52071 1548 52080
rect 162 52028 810 52037
rect 162 51994 810 52028
rect 162 51985 810 51994
rect 900 51942 1548 51951
rect 900 51908 1548 51942
rect 900 51899 1548 51908
rect 162 51856 810 51865
rect 162 51822 810 51856
rect 162 51813 810 51822
rect 900 51770 1548 51779
rect 900 51736 1548 51770
rect 900 51727 1548 51736
rect 162 51684 810 51693
rect 162 51650 810 51684
rect 162 51641 810 51650
rect 900 51598 1548 51607
rect 900 51564 1548 51598
rect 900 51555 1548 51564
rect 162 51512 810 51521
rect 162 51478 810 51512
rect 162 51469 810 51478
rect 900 51426 1548 51435
rect 900 51392 1548 51426
rect 900 51383 1548 51392
rect 162 51340 810 51349
rect 162 51306 810 51340
rect 162 51297 810 51306
rect 900 51254 1548 51263
rect 900 51220 1548 51254
rect 900 51211 1548 51220
rect 162 51168 810 51177
rect 162 51134 810 51168
rect 162 51125 810 51134
rect 900 51082 1548 51091
rect 900 51048 1548 51082
rect 900 51039 1548 51048
rect 162 50996 810 51005
rect 162 50962 810 50996
rect 162 50953 810 50962
rect 900 50910 1548 50919
rect 900 50876 1548 50910
rect 900 50867 1548 50876
rect 162 50824 810 50833
rect 162 50790 810 50824
rect 162 50781 810 50790
rect 900 50738 1548 50747
rect 900 50704 1548 50738
rect 900 50695 1548 50704
rect 162 50652 810 50661
rect 162 50618 810 50652
rect 162 50609 810 50618
rect 900 50566 1548 50575
rect 900 50532 1548 50566
rect 900 50523 1548 50532
rect 162 50480 810 50489
rect 162 50446 810 50480
rect 162 50437 810 50446
rect 900 50394 1548 50403
rect 900 50360 1548 50394
rect 900 50351 1548 50360
rect 162 50308 810 50317
rect 162 50274 810 50308
rect 162 50265 810 50274
rect 900 50222 1548 50231
rect 900 50188 1548 50222
rect 900 50179 1548 50188
rect 162 50136 810 50145
rect 162 50102 810 50136
rect 162 50093 810 50102
rect 900 50050 1548 50059
rect 900 50016 1548 50050
rect 900 50007 1548 50016
rect 162 49964 810 49973
rect 162 49930 810 49964
rect 162 49921 810 49930
rect 900 49878 1548 49887
rect 900 49844 1548 49878
rect 900 49835 1548 49844
rect 162 49792 810 49801
rect 162 49758 810 49792
rect 162 49749 810 49758
rect 900 49706 1548 49715
rect 900 49672 1548 49706
rect 900 49663 1548 49672
rect 162 49620 810 49629
rect 162 49586 810 49620
rect 162 49577 810 49586
rect 900 49534 1548 49543
rect 900 49500 1548 49534
rect 900 49491 1548 49500
rect 162 49448 810 49457
rect 162 49414 810 49448
rect 162 49405 810 49414
rect 900 49362 1548 49371
rect 900 49328 1548 49362
rect 900 49319 1548 49328
rect 162 49276 810 49285
rect 162 49242 810 49276
rect 162 49233 810 49242
rect 900 49190 1548 49199
rect 900 49156 1548 49190
rect 900 49147 1548 49156
rect 162 49104 810 49113
rect 162 49070 810 49104
rect 162 49061 810 49070
rect 900 49018 1548 49027
rect 900 48984 1548 49018
rect 900 48975 1548 48984
rect 162 48932 810 48941
rect 162 48898 810 48932
rect 162 48889 810 48898
rect 900 48846 1548 48855
rect 900 48812 1548 48846
rect 900 48803 1548 48812
rect 162 48760 810 48769
rect 162 48726 810 48760
rect 162 48717 810 48726
rect 900 48674 1548 48683
rect 900 48640 1548 48674
rect 900 48631 1548 48640
rect 162 48588 810 48597
rect 162 48554 810 48588
rect 162 48545 810 48554
rect 900 48502 1548 48511
rect 900 48468 1548 48502
rect 900 48459 1548 48468
rect 162 48416 810 48425
rect 162 48382 810 48416
rect 162 48373 810 48382
rect 900 48330 1548 48339
rect 900 48296 1548 48330
rect 900 48287 1548 48296
rect 162 48244 810 48253
rect 162 48210 810 48244
rect 162 48201 810 48210
rect 900 48158 1548 48167
rect 900 48124 1548 48158
rect 900 48115 1548 48124
rect 162 48072 810 48081
rect 162 48038 810 48072
rect 162 48029 810 48038
rect 900 47986 1548 47995
rect 900 47952 1548 47986
rect 900 47943 1548 47952
rect 162 47900 810 47909
rect 162 47866 810 47900
rect 162 47857 810 47866
rect 900 47814 1548 47823
rect 900 47780 1548 47814
rect 900 47771 1548 47780
rect 162 47728 810 47737
rect 162 47694 810 47728
rect 162 47685 810 47694
rect 900 47642 1548 47651
rect 900 47608 1548 47642
rect 900 47599 1548 47608
rect 162 47556 810 47565
rect 162 47522 810 47556
rect 162 47513 810 47522
rect 900 47470 1548 47479
rect 900 47436 1548 47470
rect 900 47427 1548 47436
rect 162 47384 810 47393
rect 162 47350 810 47384
rect 162 47341 810 47350
rect 900 47298 1548 47307
rect 900 47264 1548 47298
rect 900 47255 1548 47264
rect 162 47212 810 47221
rect 162 47178 810 47212
rect 162 47169 810 47178
rect 900 47126 1548 47135
rect 900 47092 1548 47126
rect 900 47083 1548 47092
rect 162 47040 810 47049
rect 162 47006 810 47040
rect 162 46997 810 47006
rect 900 46954 1548 46963
rect 900 46920 1548 46954
rect 900 46911 1548 46920
rect 162 46868 810 46877
rect 162 46834 810 46868
rect 162 46825 810 46834
rect 900 46782 1548 46791
rect 900 46748 1548 46782
rect 900 46739 1548 46748
rect 162 46696 810 46705
rect 162 46662 810 46696
rect 162 46653 810 46662
rect 900 46610 1548 46619
rect 900 46576 1548 46610
rect 900 46567 1548 46576
rect 162 46524 810 46533
rect 162 46490 810 46524
rect 162 46481 810 46490
rect 900 46438 1548 46447
rect 900 46404 1548 46438
rect 900 46395 1548 46404
rect 162 46352 810 46361
rect 162 46318 810 46352
rect 162 46309 810 46318
rect 900 46266 1548 46275
rect 900 46232 1548 46266
rect 900 46223 1548 46232
rect 162 46180 810 46189
rect 162 46146 810 46180
rect 162 46137 810 46146
rect 900 46094 1548 46103
rect 900 46060 1548 46094
rect 900 46051 1548 46060
rect 162 46008 810 46017
rect 162 45974 810 46008
rect 162 45965 810 45974
rect 900 45922 1548 45931
rect 900 45888 1548 45922
rect 900 45879 1548 45888
rect 162 45836 810 45845
rect 162 45802 810 45836
rect 162 45793 810 45802
rect 900 45750 1548 45759
rect 900 45716 1548 45750
rect 900 45707 1548 45716
rect 162 45664 810 45673
rect 162 45630 810 45664
rect 162 45621 810 45630
rect 900 45578 1548 45587
rect 900 45544 1548 45578
rect 900 45535 1548 45544
rect 162 45492 810 45501
rect 162 45458 810 45492
rect 162 45449 810 45458
rect 900 45406 1548 45415
rect 900 45372 1548 45406
rect 900 45363 1548 45372
rect 162 45320 810 45329
rect 162 45286 810 45320
rect 162 45277 810 45286
rect 900 45234 1548 45243
rect 900 45200 1548 45234
rect 900 45191 1548 45200
rect 162 45148 810 45157
rect 162 45114 810 45148
rect 162 45105 810 45114
rect 900 45062 1548 45071
rect 900 45028 1548 45062
rect 900 45019 1548 45028
rect 162 44976 810 44985
rect 162 44942 810 44976
rect 162 44933 810 44942
rect 900 44890 1548 44899
rect 900 44856 1548 44890
rect 900 44847 1548 44856
rect 162 44804 810 44813
rect 162 44770 810 44804
rect 162 44761 810 44770
rect 900 44718 1548 44727
rect 900 44684 1548 44718
rect 900 44675 1548 44684
rect 162 44632 810 44641
rect 162 44598 810 44632
rect 162 44589 810 44598
rect 900 44546 1548 44555
rect 900 44512 1548 44546
rect 900 44503 1548 44512
rect 162 44460 810 44469
rect 162 44426 810 44460
rect 162 44417 810 44426
rect 900 44374 1548 44383
rect 900 44340 1548 44374
rect 900 44331 1548 44340
rect 162 44288 810 44297
rect 162 44254 810 44288
rect 162 44245 810 44254
rect 900 44202 1548 44211
rect 900 44168 1548 44202
rect 900 44159 1548 44168
rect 162 44116 810 44125
rect 162 44082 810 44116
rect 162 44073 810 44082
rect 900 44030 1548 44039
rect 900 43996 1548 44030
rect 900 43987 1548 43996
rect 162 43944 810 43953
rect 162 43910 810 43944
rect 162 43901 810 43910
rect 900 43858 1548 43867
rect 900 43824 1548 43858
rect 900 43815 1548 43824
rect 162 43772 810 43781
rect 162 43738 810 43772
rect 162 43729 810 43738
rect 900 43686 1548 43695
rect 900 43652 1548 43686
rect 900 43643 1548 43652
rect 162 43600 810 43609
rect 162 43566 810 43600
rect 162 43557 810 43566
rect 900 43514 1548 43523
rect 900 43480 1548 43514
rect 900 43471 1548 43480
rect 162 43428 810 43437
rect 162 43394 810 43428
rect 162 43385 810 43394
rect 900 43342 1548 43351
rect 900 43308 1548 43342
rect 900 43299 1548 43308
rect 162 43256 810 43265
rect 162 43222 810 43256
rect 162 43213 810 43222
rect 900 43170 1548 43179
rect 900 43136 1548 43170
rect 900 43127 1548 43136
rect 162 43084 810 43093
rect 162 43050 810 43084
rect 162 43041 810 43050
rect 900 42998 1548 43007
rect 900 42964 1548 42998
rect 900 42955 1548 42964
rect 162 42912 810 42921
rect 162 42878 810 42912
rect 162 42869 810 42878
rect 900 42826 1548 42835
rect 900 42792 1548 42826
rect 900 42783 1548 42792
rect 162 42740 810 42749
rect 162 42706 810 42740
rect 162 42697 810 42706
rect 900 42654 1548 42663
rect 900 42620 1548 42654
rect 900 42611 1548 42620
rect 162 42568 810 42577
rect 162 42534 810 42568
rect 162 42525 810 42534
rect 900 42482 1548 42491
rect 900 42448 1548 42482
rect 900 42439 1548 42448
rect 162 42396 810 42405
rect 162 42362 810 42396
rect 162 42353 810 42362
rect 900 42310 1548 42319
rect 900 42276 1548 42310
rect 900 42267 1548 42276
rect 162 42224 810 42233
rect 162 42190 810 42224
rect 162 42181 810 42190
rect 900 42138 1548 42147
rect 900 42104 1548 42138
rect 900 42095 1548 42104
rect 162 42052 810 42061
rect 162 42018 810 42052
rect 162 42009 810 42018
rect 900 41966 1548 41975
rect 900 41932 1548 41966
rect 900 41923 1548 41932
rect 162 41880 810 41889
rect 162 41846 810 41880
rect 162 41837 810 41846
rect 900 41794 1548 41803
rect 900 41760 1548 41794
rect 900 41751 1548 41760
rect 162 41708 810 41717
rect 162 41674 810 41708
rect 162 41665 810 41674
rect 900 41622 1548 41631
rect 900 41588 1548 41622
rect 900 41579 1548 41588
rect 162 41536 810 41545
rect 162 41502 810 41536
rect 162 41493 810 41502
rect 900 41450 1548 41459
rect 900 41416 1548 41450
rect 900 41407 1548 41416
rect 162 41364 810 41373
rect 162 41330 810 41364
rect 162 41321 810 41330
rect 900 41278 1548 41287
rect 900 41244 1548 41278
rect 900 41235 1548 41244
rect 162 41192 810 41201
rect 162 41158 810 41192
rect 162 41149 810 41158
rect 900 41106 1548 41115
rect 900 41072 1548 41106
rect 900 41063 1548 41072
rect 162 41020 810 41029
rect 162 40986 810 41020
rect 162 40977 810 40986
rect 900 40934 1548 40943
rect 900 40900 1548 40934
rect 900 40891 1548 40900
rect 162 40848 810 40857
rect 162 40814 810 40848
rect 162 40805 810 40814
rect 900 40762 1548 40771
rect 900 40728 1548 40762
rect 900 40719 1548 40728
rect 162 40676 810 40685
rect 162 40642 810 40676
rect 162 40633 810 40642
rect 900 40590 1548 40599
rect 900 40556 1548 40590
rect 900 40547 1548 40556
rect 162 40504 810 40513
rect 162 40470 810 40504
rect 162 40461 810 40470
rect 900 40418 1548 40427
rect 900 40384 1548 40418
rect 900 40375 1548 40384
rect 162 40332 810 40341
rect 162 40298 810 40332
rect 162 40289 810 40298
rect 900 40246 1548 40255
rect 900 40212 1548 40246
rect 900 40203 1548 40212
rect 162 40160 810 40169
rect 162 40126 810 40160
rect 162 40117 810 40126
rect 900 40074 1548 40083
rect 900 40040 1548 40074
rect 900 40031 1548 40040
rect 162 39988 810 39997
rect 162 39954 810 39988
rect 162 39945 810 39954
rect 900 39902 1548 39911
rect 900 39868 1548 39902
rect 900 39859 1548 39868
rect 162 39816 810 39825
rect 162 39782 810 39816
rect 162 39773 810 39782
rect 900 39730 1548 39739
rect 900 39696 1548 39730
rect 900 39687 1548 39696
rect 162 39644 810 39653
rect 162 39610 810 39644
rect 162 39601 810 39610
rect 900 39558 1548 39567
rect 900 39524 1548 39558
rect 900 39515 1548 39524
rect 162 39472 810 39481
rect 162 39438 810 39472
rect 162 39429 810 39438
rect 900 39386 1548 39395
rect 900 39352 1548 39386
rect 900 39343 1548 39352
rect 162 39300 810 39309
rect 162 39266 810 39300
rect 162 39257 810 39266
rect 900 39214 1548 39223
rect 900 39180 1548 39214
rect 900 39171 1548 39180
rect 162 39128 810 39137
rect 162 39094 810 39128
rect 162 39085 810 39094
rect 900 39042 1548 39051
rect 900 39008 1548 39042
rect 900 38999 1548 39008
rect 162 38956 810 38965
rect 162 38922 810 38956
rect 162 38913 810 38922
rect 900 38870 1548 38879
rect 900 38836 1548 38870
rect 900 38827 1548 38836
rect 162 38784 810 38793
rect 162 38750 810 38784
rect 162 38741 810 38750
rect 900 38698 1548 38707
rect 900 38664 1548 38698
rect 900 38655 1548 38664
rect 162 38612 810 38621
rect 162 38578 810 38612
rect 162 38569 810 38578
rect 900 38526 1548 38535
rect 900 38492 1548 38526
rect 900 38483 1548 38492
rect 162 38440 810 38449
rect 162 38406 810 38440
rect 162 38397 810 38406
rect 900 38354 1548 38363
rect 900 38320 1548 38354
rect 900 38311 1548 38320
rect 162 38268 810 38277
rect 162 38234 810 38268
rect 162 38225 810 38234
rect 900 38182 1548 38191
rect 900 38148 1548 38182
rect 900 38139 1548 38148
rect 162 38096 810 38105
rect 162 38062 810 38096
rect 162 38053 810 38062
rect 900 38010 1548 38019
rect 900 37976 1548 38010
rect 900 37967 1548 37976
rect 162 37924 810 37933
rect 162 37890 810 37924
rect 162 37881 810 37890
rect 900 37838 1548 37847
rect 900 37804 1548 37838
rect 900 37795 1548 37804
rect 162 37752 810 37761
rect 162 37718 810 37752
rect 162 37709 810 37718
rect 900 37666 1548 37675
rect 900 37632 1548 37666
rect 900 37623 1548 37632
rect 162 37580 810 37589
rect 162 37546 810 37580
rect 162 37537 810 37546
rect 900 37494 1548 37503
rect 900 37460 1548 37494
rect 900 37451 1548 37460
rect 162 37408 810 37417
rect 162 37374 810 37408
rect 162 37365 810 37374
rect 900 37322 1548 37331
rect 900 37288 1548 37322
rect 900 37279 1548 37288
rect 162 37236 810 37245
rect 162 37202 810 37236
rect 162 37193 810 37202
rect 900 37150 1548 37159
rect 900 37116 1548 37150
rect 900 37107 1548 37116
rect 162 37064 810 37073
rect 162 37030 810 37064
rect 162 37021 810 37030
rect 900 36978 1548 36987
rect 900 36944 1548 36978
rect 900 36935 1548 36944
rect 162 36892 810 36901
rect 162 36858 810 36892
rect 162 36849 810 36858
rect 900 36806 1548 36815
rect 900 36772 1548 36806
rect 900 36763 1548 36772
rect 162 36720 810 36729
rect 162 36686 810 36720
rect 162 36677 810 36686
rect 900 36634 1548 36643
rect 900 36600 1548 36634
rect 900 36591 1548 36600
rect 162 36548 810 36557
rect 162 36514 810 36548
rect 162 36505 810 36514
rect 900 36462 1548 36471
rect 900 36428 1548 36462
rect 900 36419 1548 36428
rect 162 36376 810 36385
rect 162 36342 810 36376
rect 162 36333 810 36342
rect 900 36290 1548 36299
rect 900 36256 1548 36290
rect 900 36247 1548 36256
rect 162 36204 810 36213
rect 162 36170 810 36204
rect 162 36161 810 36170
rect 900 36118 1548 36127
rect 900 36084 1548 36118
rect 900 36075 1548 36084
rect 162 36032 810 36041
rect 162 35998 810 36032
rect 162 35989 810 35998
rect 900 35946 1548 35955
rect 900 35912 1548 35946
rect 900 35903 1548 35912
rect 162 35860 810 35869
rect 162 35826 810 35860
rect 162 35817 810 35826
rect 900 35774 1548 35783
rect 900 35740 1548 35774
rect 900 35731 1548 35740
rect 162 35688 810 35697
rect 162 35654 810 35688
rect 162 35645 810 35654
rect 900 35602 1548 35611
rect 900 35568 1548 35602
rect 900 35559 1548 35568
rect 162 35516 810 35525
rect 162 35482 810 35516
rect 162 35473 810 35482
rect 900 35430 1548 35439
rect 900 35396 1548 35430
rect 900 35387 1548 35396
rect 162 35344 810 35353
rect 162 35310 810 35344
rect 162 35301 810 35310
rect 900 35258 1548 35267
rect 900 35224 1548 35258
rect 900 35215 1548 35224
rect 162 35172 810 35181
rect 162 35138 810 35172
rect 162 35129 810 35138
rect 900 35086 1548 35095
rect 900 35052 1548 35086
rect 900 35043 1548 35052
rect 162 35000 810 35009
rect 162 34966 810 35000
rect 162 34957 810 34966
rect 900 34914 1548 34923
rect 900 34880 1548 34914
rect 900 34871 1548 34880
rect 162 34828 810 34837
rect 162 34794 810 34828
rect 162 34785 810 34794
rect 900 34742 1548 34751
rect 900 34708 1548 34742
rect 900 34699 1548 34708
rect 162 34656 810 34665
rect 162 34622 810 34656
rect 162 34613 810 34622
rect 900 34570 1548 34579
rect 900 34536 1548 34570
rect 900 34527 1548 34536
rect 162 34484 810 34493
rect 162 34450 810 34484
rect 162 34441 810 34450
rect 900 34398 1548 34407
rect 900 34364 1548 34398
rect 900 34355 1548 34364
rect 162 34312 810 34321
rect 162 34278 810 34312
rect 162 34269 810 34278
rect 900 34226 1548 34235
rect 900 34192 1548 34226
rect 900 34183 1548 34192
rect 162 34140 810 34149
rect 162 34106 810 34140
rect 162 34097 810 34106
rect 900 34054 1548 34063
rect 900 34020 1548 34054
rect 900 34011 1548 34020
rect 162 33968 810 33977
rect 162 33934 810 33968
rect 162 33925 810 33934
rect 900 33882 1548 33891
rect 900 33848 1548 33882
rect 900 33839 1548 33848
rect 162 33796 810 33805
rect 162 33762 810 33796
rect 162 33753 810 33762
rect 900 33710 1548 33719
rect 900 33676 1548 33710
rect 900 33667 1548 33676
rect 162 33624 810 33633
rect 162 33590 810 33624
rect 162 33581 810 33590
rect 900 33538 1548 33547
rect 900 33504 1548 33538
rect 900 33495 1548 33504
rect 162 33452 810 33461
rect 162 33418 810 33452
rect 162 33409 810 33418
rect 900 33366 1548 33375
rect 900 33332 1548 33366
rect 900 33323 1548 33332
rect 162 33280 810 33289
rect 162 33246 810 33280
rect 162 33237 810 33246
rect 900 33194 1548 33203
rect 900 33160 1548 33194
rect 900 33151 1548 33160
rect 162 33108 810 33117
rect 162 33074 810 33108
rect 162 33065 810 33074
rect 900 33022 1548 33031
rect 900 32988 1548 33022
rect 900 32979 1548 32988
rect 162 32936 810 32945
rect 162 32902 810 32936
rect 162 32893 810 32902
rect 900 32850 1548 32859
rect 900 32816 1548 32850
rect 900 32807 1548 32816
rect 162 32764 810 32773
rect 162 32730 810 32764
rect 162 32721 810 32730
rect 900 32678 1548 32687
rect 900 32644 1548 32678
rect 900 32635 1548 32644
rect 162 32592 810 32601
rect 162 32558 810 32592
rect 162 32549 810 32558
rect 900 32506 1548 32515
rect 900 32472 1548 32506
rect 900 32463 1548 32472
rect 162 32420 810 32429
rect 162 32386 810 32420
rect 162 32377 810 32386
rect 900 32334 1548 32343
rect 900 32300 1548 32334
rect 900 32291 1548 32300
rect 162 32248 810 32257
rect 162 32214 810 32248
rect 162 32205 810 32214
rect 900 32162 1548 32171
rect 900 32128 1548 32162
rect 900 32119 1548 32128
rect 162 32076 810 32085
rect 162 32042 810 32076
rect 162 32033 810 32042
rect 900 31990 1548 31999
rect 900 31956 1548 31990
rect 900 31947 1548 31956
rect 162 31904 810 31913
rect 162 31870 810 31904
rect 162 31861 810 31870
rect 900 31818 1548 31827
rect 900 31784 1548 31818
rect 900 31775 1548 31784
rect 162 31732 810 31741
rect 162 31698 810 31732
rect 162 31689 810 31698
rect 900 31646 1548 31655
rect 900 31612 1548 31646
rect 900 31603 1548 31612
rect 162 31560 810 31569
rect 162 31526 810 31560
rect 162 31517 810 31526
rect 900 31474 1548 31483
rect 900 31440 1548 31474
rect 900 31431 1548 31440
rect 162 31388 810 31397
rect 162 31354 810 31388
rect 162 31345 810 31354
rect 900 31302 1548 31311
rect 900 31268 1548 31302
rect 900 31259 1548 31268
rect 162 31216 810 31225
rect 162 31182 810 31216
rect 162 31173 810 31182
rect 900 31130 1548 31139
rect 900 31096 1548 31130
rect 900 31087 1548 31096
rect 162 31044 810 31053
rect 162 31010 810 31044
rect 162 31001 810 31010
rect 900 30958 1548 30967
rect 900 30924 1548 30958
rect 900 30915 1548 30924
rect 162 30872 810 30881
rect 162 30838 810 30872
rect 162 30829 810 30838
rect 900 30786 1548 30795
rect 900 30752 1548 30786
rect 900 30743 1548 30752
rect 162 30700 810 30709
rect 162 30666 810 30700
rect 162 30657 810 30666
rect 900 30614 1548 30623
rect 900 30580 1548 30614
rect 900 30571 1548 30580
rect 162 30528 810 30537
rect 162 30494 810 30528
rect 162 30485 810 30494
rect 900 30442 1548 30451
rect 900 30408 1548 30442
rect 900 30399 1548 30408
rect 162 30356 810 30365
rect 162 30322 810 30356
rect 162 30313 810 30322
rect 900 30270 1548 30279
rect 900 30236 1548 30270
rect 900 30227 1548 30236
rect 162 30184 810 30193
rect 162 30150 810 30184
rect 162 30141 810 30150
rect 900 30098 1548 30107
rect 900 30064 1548 30098
rect 900 30055 1548 30064
rect 162 30012 810 30021
rect 162 29978 810 30012
rect 162 29969 810 29978
rect 900 29926 1548 29935
rect 900 29892 1548 29926
rect 900 29883 1548 29892
rect 162 29840 810 29849
rect 162 29806 810 29840
rect 162 29797 810 29806
rect 900 29754 1548 29763
rect 900 29720 1548 29754
rect 900 29711 1548 29720
rect 162 29668 810 29677
rect 162 29634 810 29668
rect 162 29625 810 29634
rect 900 29582 1548 29591
rect 900 29548 1548 29582
rect 900 29539 1548 29548
rect 162 29496 810 29505
rect 162 29462 810 29496
rect 162 29453 810 29462
rect 900 29410 1548 29419
rect 900 29376 1548 29410
rect 900 29367 1548 29376
rect 162 29324 810 29333
rect 162 29290 810 29324
rect 162 29281 810 29290
rect 900 29238 1548 29247
rect 900 29204 1548 29238
rect 900 29195 1548 29204
rect 162 29152 810 29161
rect 162 29118 810 29152
rect 162 29109 810 29118
rect 900 29066 1548 29075
rect 900 29032 1548 29066
rect 900 29023 1548 29032
rect 162 28980 810 28989
rect 162 28946 810 28980
rect 162 28937 810 28946
rect 900 28894 1548 28903
rect 900 28860 1548 28894
rect 900 28851 1548 28860
rect 162 28808 810 28817
rect 162 28774 810 28808
rect 162 28765 810 28774
rect 900 28722 1548 28731
rect 900 28688 1548 28722
rect 900 28679 1548 28688
rect 162 28636 810 28645
rect 162 28602 810 28636
rect 162 28593 810 28602
rect 900 28550 1548 28559
rect 900 28516 1548 28550
rect 900 28507 1548 28516
rect 162 28464 810 28473
rect 162 28430 810 28464
rect 162 28421 810 28430
rect 900 28378 1548 28387
rect 900 28344 1548 28378
rect 900 28335 1548 28344
rect 162 28292 810 28301
rect 162 28258 810 28292
rect 162 28249 810 28258
rect 900 28206 1548 28215
rect 900 28172 1548 28206
rect 900 28163 1548 28172
rect 162 28120 810 28129
rect 162 28086 810 28120
rect 162 28077 810 28086
rect 900 28034 1548 28043
rect 900 28000 1548 28034
rect 900 27991 1548 28000
rect 162 27948 810 27957
rect 162 27914 810 27948
rect 162 27905 810 27914
rect 900 27862 1548 27871
rect 900 27828 1548 27862
rect 900 27819 1548 27828
rect 162 27776 810 27785
rect 162 27742 810 27776
rect 162 27733 810 27742
rect 900 27690 1548 27699
rect 900 27656 1548 27690
rect 900 27647 1548 27656
rect 162 27604 810 27613
rect 162 27570 810 27604
rect 162 27561 810 27570
rect 900 27518 1548 27527
rect 900 27484 1548 27518
rect 900 27475 1548 27484
rect 162 27432 810 27441
rect 162 27398 810 27432
rect 162 27389 810 27398
rect 900 27346 1548 27355
rect 900 27312 1548 27346
rect 900 27303 1548 27312
rect 162 27260 810 27269
rect 162 27226 810 27260
rect 162 27217 810 27226
rect 900 27174 1548 27183
rect 900 27140 1548 27174
rect 900 27131 1548 27140
rect 162 27088 810 27097
rect 162 27054 810 27088
rect 162 27045 810 27054
rect 900 27002 1548 27011
rect 900 26968 1548 27002
rect 900 26959 1548 26968
rect 162 26916 810 26925
rect 162 26882 810 26916
rect 162 26873 810 26882
rect 900 26830 1548 26839
rect 900 26796 1548 26830
rect 900 26787 1548 26796
rect 162 26744 810 26753
rect 162 26710 810 26744
rect 162 26701 810 26710
rect 900 26658 1548 26667
rect 900 26624 1548 26658
rect 900 26615 1548 26624
rect 162 26572 810 26581
rect 162 26538 810 26572
rect 162 26529 810 26538
rect 900 26486 1548 26495
rect 900 26452 1548 26486
rect 900 26443 1548 26452
rect 162 26400 810 26409
rect 162 26366 810 26400
rect 162 26357 810 26366
rect 900 26314 1548 26323
rect 900 26280 1548 26314
rect 900 26271 1548 26280
rect 162 26228 810 26237
rect 162 26194 810 26228
rect 162 26185 810 26194
rect 900 26142 1548 26151
rect 900 26108 1548 26142
rect 900 26099 1548 26108
rect 162 26056 810 26065
rect 162 26022 810 26056
rect 162 26013 810 26022
rect 900 25970 1548 25979
rect 900 25936 1548 25970
rect 900 25927 1548 25936
rect 162 25884 810 25893
rect 162 25850 810 25884
rect 162 25841 810 25850
rect 900 25798 1548 25807
rect 900 25764 1548 25798
rect 900 25755 1548 25764
rect 162 25712 810 25721
rect 162 25678 810 25712
rect 162 25669 810 25678
rect 900 25626 1548 25635
rect 900 25592 1548 25626
rect 900 25583 1548 25592
rect 162 25540 810 25549
rect 162 25506 810 25540
rect 162 25497 810 25506
rect 900 25454 1548 25463
rect 900 25420 1548 25454
rect 900 25411 1548 25420
rect 162 25368 810 25377
rect 162 25334 810 25368
rect 162 25325 810 25334
rect 900 25282 1548 25291
rect 900 25248 1548 25282
rect 900 25239 1548 25248
rect 162 25196 810 25205
rect 162 25162 810 25196
rect 162 25153 810 25162
rect 900 25110 1548 25119
rect 900 25076 1548 25110
rect 900 25067 1548 25076
rect 162 25024 810 25033
rect 162 24990 810 25024
rect 162 24981 810 24990
rect 900 24938 1548 24947
rect 900 24904 1548 24938
rect 900 24895 1548 24904
rect 162 24852 810 24861
rect 162 24818 810 24852
rect 162 24809 810 24818
rect 900 24766 1548 24775
rect 900 24732 1548 24766
rect 900 24723 1548 24732
rect 162 24680 810 24689
rect 162 24646 810 24680
rect 162 24637 810 24646
rect 900 24594 1548 24603
rect 900 24560 1548 24594
rect 900 24551 1548 24560
rect 162 24508 810 24517
rect 162 24474 810 24508
rect 162 24465 810 24474
rect 900 24422 1548 24431
rect 900 24388 1548 24422
rect 900 24379 1548 24388
rect 162 24336 810 24345
rect 162 24302 810 24336
rect 162 24293 810 24302
rect 900 24250 1548 24259
rect 900 24216 1548 24250
rect 900 24207 1548 24216
rect 162 24164 810 24173
rect 162 24130 810 24164
rect 162 24121 810 24130
rect 900 24078 1548 24087
rect 900 24044 1548 24078
rect 900 24035 1548 24044
rect 162 23992 810 24001
rect 162 23958 810 23992
rect 162 23949 810 23958
rect 900 23906 1548 23915
rect 900 23872 1548 23906
rect 900 23863 1548 23872
rect 162 23820 810 23829
rect 162 23786 810 23820
rect 162 23777 810 23786
rect 900 23734 1548 23743
rect 900 23700 1548 23734
rect 900 23691 1548 23700
rect 162 23648 810 23657
rect 162 23614 810 23648
rect 162 23605 810 23614
rect 900 23562 1548 23571
rect 900 23528 1548 23562
rect 900 23519 1548 23528
rect 162 23476 810 23485
rect 162 23442 810 23476
rect 162 23433 810 23442
rect 900 23390 1548 23399
rect 900 23356 1548 23390
rect 900 23347 1548 23356
rect 162 23304 810 23313
rect 162 23270 810 23304
rect 162 23261 810 23270
rect 900 23218 1548 23227
rect 900 23184 1548 23218
rect 900 23175 1548 23184
rect 162 23132 810 23141
rect 162 23098 810 23132
rect 162 23089 810 23098
rect 900 23046 1548 23055
rect 900 23012 1548 23046
rect 900 23003 1548 23012
rect 162 22960 810 22969
rect 162 22926 810 22960
rect 162 22917 810 22926
rect 900 22874 1548 22883
rect 900 22840 1548 22874
rect 900 22831 1548 22840
rect 162 22788 810 22797
rect 162 22754 810 22788
rect 162 22745 810 22754
rect 900 22702 1548 22711
rect 900 22668 1548 22702
rect 900 22659 1548 22668
rect 162 22616 810 22625
rect 162 22582 810 22616
rect 162 22573 810 22582
rect 900 22530 1548 22539
rect 900 22496 1548 22530
rect 900 22487 1548 22496
rect 162 22444 810 22453
rect 162 22410 810 22444
rect 162 22401 810 22410
rect 900 22358 1548 22367
rect 900 22324 1548 22358
rect 900 22315 1548 22324
rect 162 22272 810 22281
rect 162 22238 810 22272
rect 162 22229 810 22238
rect 900 22186 1548 22195
rect 900 22152 1548 22186
rect 900 22143 1548 22152
rect 162 22100 810 22109
rect 162 22066 810 22100
rect 162 22057 810 22066
rect 900 22014 1548 22023
rect 900 21980 1548 22014
rect 900 21971 1548 21980
rect 162 21928 810 21937
rect 162 21894 810 21928
rect 162 21885 810 21894
rect 900 21842 1548 21851
rect 900 21808 1548 21842
rect 900 21799 1548 21808
rect 162 21756 810 21765
rect 162 21722 810 21756
rect 162 21713 810 21722
rect 900 21670 1548 21679
rect 900 21636 1548 21670
rect 900 21627 1548 21636
rect 162 21584 810 21593
rect 162 21550 810 21584
rect 162 21541 810 21550
rect 900 21498 1548 21507
rect 900 21464 1548 21498
rect 900 21455 1548 21464
rect 162 21412 810 21421
rect 162 21378 810 21412
rect 162 21369 810 21378
rect 900 21326 1548 21335
rect 900 21292 1548 21326
rect 900 21283 1548 21292
rect 162 21240 810 21249
rect 162 21206 810 21240
rect 162 21197 810 21206
rect 900 21154 1548 21163
rect 900 21120 1548 21154
rect 900 21111 1548 21120
rect 162 21068 810 21077
rect 162 21034 810 21068
rect 162 21025 810 21034
rect 900 20982 1548 20991
rect 900 20948 1548 20982
rect 900 20939 1548 20948
rect 162 20896 810 20905
rect 162 20862 810 20896
rect 162 20853 810 20862
rect 900 20810 1548 20819
rect 900 20776 1548 20810
rect 900 20767 1548 20776
rect 162 20724 810 20733
rect 162 20690 810 20724
rect 162 20681 810 20690
rect 900 20638 1548 20647
rect 900 20604 1548 20638
rect 900 20595 1548 20604
rect 162 20552 810 20561
rect 162 20518 810 20552
rect 162 20509 810 20518
rect 900 20466 1548 20475
rect 900 20432 1548 20466
rect 900 20423 1548 20432
rect 162 20380 810 20389
rect 162 20346 810 20380
rect 162 20337 810 20346
rect 900 20294 1548 20303
rect 900 20260 1548 20294
rect 900 20251 1548 20260
rect 162 20208 810 20217
rect 162 20174 810 20208
rect 162 20165 810 20174
rect 900 20122 1548 20131
rect 900 20088 1548 20122
rect 900 20079 1548 20088
rect 162 20036 810 20045
rect 162 20002 810 20036
rect 162 19993 810 20002
rect 900 19950 1548 19959
rect 900 19916 1548 19950
rect 900 19907 1548 19916
rect 162 19864 810 19873
rect 162 19830 810 19864
rect 162 19821 810 19830
rect 900 19778 1548 19787
rect 900 19744 1548 19778
rect 900 19735 1548 19744
rect 162 19692 810 19701
rect 162 19658 810 19692
rect 162 19649 810 19658
rect 900 19606 1548 19615
rect 900 19572 1548 19606
rect 900 19563 1548 19572
rect 162 19520 810 19529
rect 162 19486 810 19520
rect 162 19477 810 19486
rect 900 19434 1548 19443
rect 900 19400 1548 19434
rect 900 19391 1548 19400
rect 162 19348 810 19357
rect 162 19314 810 19348
rect 162 19305 810 19314
rect 900 19262 1548 19271
rect 900 19228 1548 19262
rect 900 19219 1548 19228
rect 162 19176 810 19185
rect 162 19142 810 19176
rect 162 19133 810 19142
rect 900 19090 1548 19099
rect 900 19056 1548 19090
rect 900 19047 1548 19056
rect 162 19004 810 19013
rect 162 18970 810 19004
rect 162 18961 810 18970
rect 900 18918 1548 18927
rect 900 18884 1548 18918
rect 900 18875 1548 18884
rect 162 18832 810 18841
rect 162 18798 810 18832
rect 162 18789 810 18798
rect 900 18746 1548 18755
rect 900 18712 1548 18746
rect 900 18703 1548 18712
rect 162 18660 810 18669
rect 162 18626 810 18660
rect 162 18617 810 18626
rect 900 18574 1548 18583
rect 900 18540 1548 18574
rect 900 18531 1548 18540
rect 162 18488 810 18497
rect 162 18454 810 18488
rect 162 18445 810 18454
rect 900 18402 1548 18411
rect 900 18368 1548 18402
rect 900 18359 1548 18368
rect 162 18316 810 18325
rect 162 18282 810 18316
rect 162 18273 810 18282
rect 900 18230 1548 18239
rect 900 18196 1548 18230
rect 900 18187 1548 18196
rect 162 18144 810 18153
rect 162 18110 810 18144
rect 162 18101 810 18110
rect 900 18058 1548 18067
rect 900 18024 1548 18058
rect 900 18015 1548 18024
rect 162 17972 810 17981
rect 162 17938 810 17972
rect 162 17929 810 17938
rect 900 17886 1548 17895
rect 900 17852 1548 17886
rect 900 17843 1548 17852
rect 162 17800 810 17809
rect 162 17766 810 17800
rect 162 17757 810 17766
rect 900 17714 1548 17723
rect 900 17680 1548 17714
rect 900 17671 1548 17680
rect 162 17628 810 17637
rect 162 17594 810 17628
rect 162 17585 810 17594
rect 900 17542 1548 17551
rect 900 17508 1548 17542
rect 900 17499 1548 17508
rect 162 17456 810 17465
rect 162 17422 810 17456
rect 162 17413 810 17422
rect 900 17370 1548 17379
rect 900 17336 1548 17370
rect 900 17327 1548 17336
rect 162 17284 810 17293
rect 162 17250 810 17284
rect 162 17241 810 17250
rect 900 17198 1548 17207
rect 900 17164 1548 17198
rect 900 17155 1548 17164
rect 162 17112 810 17121
rect 162 17078 810 17112
rect 162 17069 810 17078
rect 900 17026 1548 17035
rect 900 16992 1548 17026
rect 900 16983 1548 16992
rect 162 16940 810 16949
rect 162 16906 810 16940
rect 162 16897 810 16906
rect 900 16854 1548 16863
rect 900 16820 1548 16854
rect 900 16811 1548 16820
rect 162 16768 810 16777
rect 162 16734 810 16768
rect 162 16725 810 16734
rect 900 16682 1548 16691
rect 900 16648 1548 16682
rect 900 16639 1548 16648
rect 162 16596 810 16605
rect 162 16562 810 16596
rect 162 16553 810 16562
rect 900 16510 1548 16519
rect 900 16476 1548 16510
rect 900 16467 1548 16476
rect 162 16424 810 16433
rect 162 16390 810 16424
rect 162 16381 810 16390
rect 900 16338 1548 16347
rect 900 16304 1548 16338
rect 900 16295 1548 16304
rect 162 16252 810 16261
rect 162 16218 810 16252
rect 162 16209 810 16218
rect 900 16166 1548 16175
rect 900 16132 1548 16166
rect 900 16123 1548 16132
rect 162 16080 810 16089
rect 162 16046 810 16080
rect 162 16037 810 16046
rect 900 15994 1548 16003
rect 900 15960 1548 15994
rect 900 15951 1548 15960
rect 162 15908 810 15917
rect 162 15874 810 15908
rect 162 15865 810 15874
rect 900 15822 1548 15831
rect 900 15788 1548 15822
rect 900 15779 1548 15788
rect 162 15736 810 15745
rect 162 15702 810 15736
rect 162 15693 810 15702
rect 900 15650 1548 15659
rect 900 15616 1548 15650
rect 900 15607 1548 15616
rect 162 15564 810 15573
rect 162 15530 810 15564
rect 162 15521 810 15530
rect 900 15478 1548 15487
rect 900 15444 1548 15478
rect 900 15435 1548 15444
rect 162 15392 810 15401
rect 162 15358 810 15392
rect 162 15349 810 15358
rect 900 15306 1548 15315
rect 900 15272 1548 15306
rect 900 15263 1548 15272
rect 162 15220 810 15229
rect 162 15186 810 15220
rect 162 15177 810 15186
rect 900 15134 1548 15143
rect 900 15100 1548 15134
rect 900 15091 1548 15100
rect 162 15048 810 15057
rect 162 15014 810 15048
rect 162 15005 810 15014
rect 900 14962 1548 14971
rect 900 14928 1548 14962
rect 900 14919 1548 14928
rect 162 14876 810 14885
rect 162 14842 810 14876
rect 162 14833 810 14842
rect 900 14790 1548 14799
rect 900 14756 1548 14790
rect 900 14747 1548 14756
rect 162 14704 810 14713
rect 162 14670 810 14704
rect 162 14661 810 14670
rect 900 14618 1548 14627
rect 900 14584 1548 14618
rect 900 14575 1548 14584
rect 162 14532 810 14541
rect 162 14498 810 14532
rect 162 14489 810 14498
rect 900 14446 1548 14455
rect 900 14412 1548 14446
rect 900 14403 1548 14412
rect 162 14360 810 14369
rect 162 14326 810 14360
rect 162 14317 810 14326
rect 900 14274 1548 14283
rect 900 14240 1548 14274
rect 900 14231 1548 14240
rect 162 14188 810 14197
rect 162 14154 810 14188
rect 162 14145 810 14154
rect 900 14102 1548 14111
rect 900 14068 1548 14102
rect 900 14059 1548 14068
rect 162 14016 810 14025
rect 162 13982 810 14016
rect 162 13973 810 13982
rect 900 13930 1548 13939
rect 900 13896 1548 13930
rect 900 13887 1548 13896
rect 162 13844 810 13853
rect 162 13810 810 13844
rect 162 13801 810 13810
rect 900 13758 1548 13767
rect 900 13724 1548 13758
rect 900 13715 1548 13724
rect 162 13672 810 13681
rect 162 13638 810 13672
rect 162 13629 810 13638
rect 900 13586 1548 13595
rect 900 13552 1548 13586
rect 900 13543 1548 13552
rect 162 13500 810 13509
rect 162 13466 810 13500
rect 162 13457 810 13466
rect 900 13414 1548 13423
rect 900 13380 1548 13414
rect 900 13371 1548 13380
rect 162 13328 810 13337
rect 162 13294 810 13328
rect 162 13285 810 13294
rect 900 13242 1548 13251
rect 900 13208 1548 13242
rect 900 13199 1548 13208
rect 162 13156 810 13165
rect 162 13122 810 13156
rect 162 13113 810 13122
rect 900 13070 1548 13079
rect 900 13036 1548 13070
rect 900 13027 1548 13036
rect 162 12984 810 12993
rect 162 12950 810 12984
rect 162 12941 810 12950
rect 900 12898 1548 12907
rect 900 12864 1548 12898
rect 900 12855 1548 12864
rect 162 12812 810 12821
rect 162 12778 810 12812
rect 162 12769 810 12778
rect 900 12726 1548 12735
rect 900 12692 1548 12726
rect 900 12683 1548 12692
rect 162 12640 810 12649
rect 162 12606 810 12640
rect 162 12597 810 12606
rect 900 12554 1548 12563
rect 900 12520 1548 12554
rect 900 12511 1548 12520
rect 162 12468 810 12477
rect 162 12434 810 12468
rect 162 12425 810 12434
rect 900 12382 1548 12391
rect 900 12348 1548 12382
rect 900 12339 1548 12348
rect 162 12296 810 12305
rect 162 12262 810 12296
rect 162 12253 810 12262
rect 900 12210 1548 12219
rect 900 12176 1548 12210
rect 900 12167 1548 12176
rect 162 12124 810 12133
rect 162 12090 810 12124
rect 162 12081 810 12090
rect 900 12038 1548 12047
rect 900 12004 1548 12038
rect 900 11995 1548 12004
rect 162 11952 810 11961
rect 162 11918 810 11952
rect 162 11909 810 11918
rect 900 11866 1548 11875
rect 900 11832 1548 11866
rect 900 11823 1548 11832
rect 162 11780 810 11789
rect 162 11746 810 11780
rect 162 11737 810 11746
rect 900 11694 1548 11703
rect 900 11660 1548 11694
rect 900 11651 1548 11660
rect 162 11608 810 11617
rect 162 11574 810 11608
rect 162 11565 810 11574
rect 900 11522 1548 11531
rect 900 11488 1548 11522
rect 900 11479 1548 11488
rect 162 11436 810 11445
rect 162 11402 810 11436
rect 162 11393 810 11402
rect 900 11350 1548 11359
rect 900 11316 1548 11350
rect 900 11307 1548 11316
rect 162 11264 810 11273
rect 162 11230 810 11264
rect 162 11221 810 11230
rect 900 11178 1548 11187
rect 900 11144 1548 11178
rect 900 11135 1548 11144
rect 162 11092 810 11101
rect 162 11058 810 11092
rect 162 11049 810 11058
rect 900 11006 1548 11015
rect 900 10972 1548 11006
rect 900 10963 1548 10972
rect 162 10920 810 10929
rect 162 10886 810 10920
rect 162 10877 810 10886
rect 900 10834 1548 10843
rect 900 10800 1548 10834
rect 900 10791 1548 10800
rect 162 10748 810 10757
rect 162 10714 810 10748
rect 162 10705 810 10714
rect 900 10662 1548 10671
rect 900 10628 1548 10662
rect 900 10619 1548 10628
rect 162 10576 810 10585
rect 162 10542 810 10576
rect 162 10533 810 10542
rect 900 10490 1548 10499
rect 900 10456 1548 10490
rect 900 10447 1548 10456
rect 162 10404 810 10413
rect 162 10370 810 10404
rect 162 10361 810 10370
rect 900 10318 1548 10327
rect 900 10284 1548 10318
rect 900 10275 1548 10284
rect 162 10232 810 10241
rect 162 10198 810 10232
rect 162 10189 810 10198
rect 900 10146 1548 10155
rect 900 10112 1548 10146
rect 900 10103 1548 10112
rect 162 10060 810 10069
rect 162 10026 810 10060
rect 162 10017 810 10026
rect 900 9974 1548 9983
rect 900 9940 1548 9974
rect 900 9931 1548 9940
rect 162 9888 810 9897
rect 162 9854 810 9888
rect 162 9845 810 9854
rect 900 9802 1548 9811
rect 900 9768 1548 9802
rect 900 9759 1548 9768
rect 162 9716 810 9725
rect 162 9682 810 9716
rect 162 9673 810 9682
rect 900 9630 1548 9639
rect 900 9596 1548 9630
rect 900 9587 1548 9596
rect 162 9544 810 9553
rect 162 9510 810 9544
rect 162 9501 810 9510
rect 900 9458 1548 9467
rect 900 9424 1548 9458
rect 900 9415 1548 9424
rect 162 9372 810 9381
rect 162 9338 810 9372
rect 162 9329 810 9338
rect 900 9286 1548 9295
rect 900 9252 1548 9286
rect 900 9243 1548 9252
rect 162 9200 810 9209
rect 162 9166 810 9200
rect 162 9157 810 9166
rect 900 9114 1548 9123
rect 900 9080 1548 9114
rect 900 9071 1548 9080
rect 162 9028 810 9037
rect 162 8994 810 9028
rect 162 8985 810 8994
rect 900 8942 1548 8951
rect 900 8908 1548 8942
rect 900 8899 1548 8908
rect 162 8856 810 8865
rect 162 8822 810 8856
rect 162 8813 810 8822
rect 900 8770 1548 8779
rect 900 8736 1548 8770
rect 900 8727 1548 8736
rect 162 8684 810 8693
rect 162 8650 810 8684
rect 162 8641 810 8650
rect 900 8598 1548 8607
rect 900 8564 1548 8598
rect 900 8555 1548 8564
rect 162 8512 810 8521
rect 162 8478 810 8512
rect 162 8469 810 8478
rect 900 8426 1548 8435
rect 900 8392 1548 8426
rect 900 8383 1548 8392
rect 162 8340 810 8349
rect 162 8306 810 8340
rect 162 8297 810 8306
rect 900 8254 1548 8263
rect 900 8220 1548 8254
rect 900 8211 1548 8220
rect 162 8168 810 8177
rect 162 8134 810 8168
rect 162 8125 810 8134
rect 900 8082 1548 8091
rect 900 8048 1548 8082
rect 900 8039 1548 8048
rect 162 7996 810 8005
rect 162 7962 810 7996
rect 162 7953 810 7962
rect 900 7910 1548 7919
rect 900 7876 1548 7910
rect 900 7867 1548 7876
rect 162 7824 810 7833
rect 162 7790 810 7824
rect 162 7781 810 7790
rect 900 7738 1548 7747
rect 900 7704 1548 7738
rect 900 7695 1548 7704
rect 162 7652 810 7661
rect 162 7618 810 7652
rect 162 7609 810 7618
rect 900 7566 1548 7575
rect 900 7532 1548 7566
rect 900 7523 1548 7532
rect 162 7480 810 7489
rect 162 7446 810 7480
rect 162 7437 810 7446
rect 900 7394 1548 7403
rect 900 7360 1548 7394
rect 900 7351 1548 7360
rect 162 7308 810 7317
rect 162 7274 810 7308
rect 162 7265 810 7274
rect 900 7222 1548 7231
rect 900 7188 1548 7222
rect 900 7179 1548 7188
rect 162 7136 810 7145
rect 162 7102 810 7136
rect 162 7093 810 7102
rect 900 7050 1548 7059
rect 900 7016 1548 7050
rect 900 7007 1548 7016
rect 162 6964 810 6973
rect 162 6930 810 6964
rect 162 6921 810 6930
rect 900 6878 1548 6887
rect 900 6844 1548 6878
rect 900 6835 1548 6844
rect 162 6792 810 6801
rect 162 6758 810 6792
rect 162 6749 810 6758
rect 900 6706 1548 6715
rect 900 6672 1548 6706
rect 900 6663 1548 6672
rect 162 6620 810 6629
rect 162 6586 810 6620
rect 162 6577 810 6586
rect 900 6534 1548 6543
rect 900 6500 1548 6534
rect 900 6491 1548 6500
rect 162 6448 810 6457
rect 162 6414 810 6448
rect 162 6405 810 6414
rect 900 6362 1548 6371
rect 900 6328 1548 6362
rect 900 6319 1548 6328
rect 162 6276 810 6285
rect 162 6242 810 6276
rect 162 6233 810 6242
rect 900 6190 1548 6199
rect 900 6156 1548 6190
rect 900 6147 1548 6156
rect 162 6104 810 6113
rect 162 6070 810 6104
rect 162 6061 810 6070
rect 900 6018 1548 6027
rect 900 5984 1548 6018
rect 900 5975 1548 5984
rect 162 5932 810 5941
rect 162 5898 810 5932
rect 162 5889 810 5898
rect 900 5846 1548 5855
rect 900 5812 1548 5846
rect 900 5803 1548 5812
rect 162 5760 810 5769
rect 162 5726 810 5760
rect 162 5717 810 5726
rect 900 5674 1548 5683
rect 900 5640 1548 5674
rect 900 5631 1548 5640
rect 162 5588 810 5597
rect 162 5554 810 5588
rect 162 5545 810 5554
rect 900 5502 1548 5511
rect 900 5468 1548 5502
rect 900 5459 1548 5468
rect 162 5416 810 5425
rect 162 5382 810 5416
rect 162 5373 810 5382
rect 900 5330 1548 5339
rect 900 5296 1548 5330
rect 900 5287 1548 5296
rect 162 5244 810 5253
rect 162 5210 810 5244
rect 162 5201 810 5210
rect 900 5158 1548 5167
rect 900 5124 1548 5158
rect 900 5115 1548 5124
rect 162 5072 810 5081
rect 162 5038 810 5072
rect 162 5029 810 5038
rect 900 4986 1548 4995
rect 900 4952 1548 4986
rect 900 4943 1548 4952
rect 162 4900 810 4909
rect 162 4866 810 4900
rect 162 4857 810 4866
rect 900 4814 1548 4823
rect 900 4780 1548 4814
rect 900 4771 1548 4780
rect 162 4728 810 4737
rect 162 4694 810 4728
rect 162 4685 810 4694
rect 900 4642 1548 4651
rect 900 4608 1548 4642
rect 900 4599 1548 4608
rect 162 4556 810 4565
rect 162 4522 810 4556
rect 162 4513 810 4522
rect 900 4470 1548 4479
rect 900 4436 1548 4470
rect 900 4427 1548 4436
rect 162 4384 810 4393
rect 162 4350 810 4384
rect 162 4341 810 4350
rect 900 4298 1548 4307
rect 900 4264 1548 4298
rect 900 4255 1548 4264
rect 162 4212 810 4221
rect 162 4178 810 4212
rect 162 4169 810 4178
rect 900 4126 1548 4135
rect 900 4092 1548 4126
rect 900 4083 1548 4092
rect 162 4040 810 4049
rect 162 4006 810 4040
rect 162 3997 810 4006
rect 900 3954 1548 3963
rect 900 3920 1548 3954
rect 900 3911 1548 3920
rect 162 3868 810 3877
rect 162 3834 810 3868
rect 162 3825 810 3834
rect 900 3782 1548 3791
rect 900 3748 1548 3782
rect 900 3739 1548 3748
rect 162 3696 810 3705
rect 162 3662 810 3696
rect 162 3653 810 3662
rect 900 3610 1548 3619
rect 900 3576 1548 3610
rect 900 3567 1548 3576
rect 162 3524 810 3533
rect 162 3490 810 3524
rect 162 3481 810 3490
rect 900 3438 1548 3447
rect 900 3404 1548 3438
rect 900 3395 1548 3404
rect 162 3352 810 3361
rect 162 3318 810 3352
rect 162 3309 810 3318
rect 900 3266 1548 3275
rect 900 3232 1548 3266
rect 900 3223 1548 3232
rect 162 3180 810 3189
rect 162 3146 810 3180
rect 162 3137 810 3146
rect 900 3094 1548 3103
rect 900 3060 1548 3094
rect 900 3051 1548 3060
rect 162 3008 810 3017
rect 162 2974 810 3008
rect 162 2965 810 2974
rect 900 2922 1548 2931
rect 900 2888 1548 2922
rect 900 2879 1548 2888
rect 162 2836 810 2845
rect 162 2802 810 2836
rect 162 2793 810 2802
rect 900 2750 1548 2759
rect 900 2716 1548 2750
rect 900 2707 1548 2716
rect 162 2664 810 2673
rect 162 2630 810 2664
rect 162 2621 810 2630
rect 900 2578 1548 2587
rect 900 2544 1548 2578
rect 900 2535 1548 2544
rect 162 2492 810 2501
rect 162 2458 810 2492
rect 162 2449 810 2458
rect 900 2406 1548 2415
rect 900 2372 1548 2406
rect 900 2363 1548 2372
rect 162 2320 810 2329
rect 162 2286 810 2320
rect 162 2277 810 2286
rect 900 2234 1548 2243
rect 900 2200 1548 2234
rect 900 2191 1548 2200
rect 162 2148 810 2157
rect 162 2114 810 2148
rect 162 2105 810 2114
rect 900 2062 1548 2071
rect 900 2028 1548 2062
rect 900 2019 1548 2028
rect 162 1976 810 1985
rect 162 1942 810 1976
rect 162 1933 810 1942
rect 900 1890 1548 1899
rect 900 1856 1548 1890
rect 900 1847 1548 1856
rect 162 1804 810 1813
rect 162 1770 810 1804
rect 162 1761 810 1770
rect 900 1718 1548 1727
rect 900 1684 1548 1718
rect 900 1675 1548 1684
rect 162 1632 810 1641
rect 162 1598 810 1632
rect 162 1589 810 1598
rect 900 1546 1548 1555
rect 900 1512 1548 1546
rect 900 1503 1548 1512
rect 162 1460 810 1469
rect 162 1426 810 1460
rect 162 1417 810 1426
rect 900 1374 1548 1383
rect 900 1340 1548 1374
rect 900 1331 1548 1340
rect 162 1288 810 1297
rect 162 1254 810 1288
rect 162 1245 810 1254
rect 900 1202 1548 1211
rect 900 1168 1548 1202
rect 900 1159 1548 1168
rect 162 1116 810 1125
rect 162 1082 810 1116
rect 162 1073 810 1082
rect 900 1030 1548 1039
rect 900 996 1548 1030
rect 900 987 1548 996
rect 162 944 810 953
rect 162 910 810 944
rect 162 901 810 910
rect 900 858 1548 867
rect 900 824 1548 858
rect 900 815 1548 824
rect 162 772 810 781
rect 162 738 810 772
rect 162 729 810 738
rect 900 686 1548 695
rect 900 652 1548 686
rect 900 643 1548 652
rect 162 600 810 609
rect 162 566 810 600
rect 162 557 810 566
rect 900 514 1548 523
rect 900 480 1548 514
rect 900 471 1548 480
rect 162 428 810 437
rect 162 394 810 428
rect 162 385 810 394
rect 900 342 1548 351
rect 900 308 1548 342
rect 900 299 1548 308
rect 162 256 810 265
rect 162 222 810 256
rect 162 213 810 222
rect 1618 179 1628 100059
rect 1628 179 1662 100059
rect 1662 179 1672 100059
rect 900 170 1548 179
rect 900 136 1548 170
rect 1618 169 1672 179
rect 900 127 1548 136
<< metal2 >>
rect 156 100025 816 100111
rect 156 99973 162 100025
rect 810 99973 816 100025
rect 156 99853 816 99973
rect 156 99801 162 99853
rect 810 99801 816 99853
rect 156 99681 816 99801
rect 156 99629 162 99681
rect 810 99629 816 99681
rect 156 99509 816 99629
rect 156 99457 162 99509
rect 810 99457 816 99509
rect 156 99337 816 99457
rect 156 99285 162 99337
rect 810 99285 816 99337
rect 156 99165 816 99285
rect 156 99113 162 99165
rect 810 99113 816 99165
rect 156 98993 816 99113
rect 156 98941 162 98993
rect 810 98941 816 98993
rect 156 98821 816 98941
rect 156 98769 162 98821
rect 810 98769 816 98821
rect 156 98649 816 98769
rect 156 98597 162 98649
rect 810 98597 816 98649
rect 156 98477 816 98597
rect 156 98425 162 98477
rect 810 98425 816 98477
rect 156 98305 816 98425
rect 156 98253 162 98305
rect 810 98253 816 98305
rect 156 98133 816 98253
rect 156 98081 162 98133
rect 810 98081 816 98133
rect 156 97961 816 98081
rect 156 97909 162 97961
rect 810 97909 816 97961
rect 156 97789 816 97909
rect 156 97737 162 97789
rect 810 97737 816 97789
rect 156 97617 816 97737
rect 156 97565 162 97617
rect 810 97565 816 97617
rect 156 97445 816 97565
rect 156 97393 162 97445
rect 810 97393 816 97445
rect 156 97273 816 97393
rect 156 97221 162 97273
rect 810 97221 816 97273
rect 156 97101 816 97221
rect 156 97049 162 97101
rect 810 97049 816 97101
rect 156 96929 816 97049
rect 156 96877 162 96929
rect 810 96877 816 96929
rect 156 96757 816 96877
rect 156 96705 162 96757
rect 810 96705 816 96757
rect 156 96585 816 96705
rect 156 96533 162 96585
rect 810 96533 816 96585
rect 156 96413 816 96533
rect 156 96361 162 96413
rect 810 96361 816 96413
rect 156 96241 816 96361
rect 156 96189 162 96241
rect 810 96189 816 96241
rect 156 96069 816 96189
rect 156 96017 162 96069
rect 810 96017 816 96069
rect 156 95897 816 96017
rect 156 95845 162 95897
rect 810 95845 816 95897
rect 156 95725 816 95845
rect 156 95673 162 95725
rect 810 95673 816 95725
rect 156 95553 816 95673
rect 156 95501 162 95553
rect 810 95501 816 95553
rect 156 95381 816 95501
rect 156 95329 162 95381
rect 810 95329 816 95381
rect 156 95209 816 95329
rect 156 95157 162 95209
rect 810 95157 816 95209
rect 156 95037 816 95157
rect 156 94985 162 95037
rect 810 94985 816 95037
rect 156 94865 816 94985
rect 156 94813 162 94865
rect 810 94813 816 94865
rect 156 94693 816 94813
rect 156 94641 162 94693
rect 810 94641 816 94693
rect 156 94521 816 94641
rect 156 94469 162 94521
rect 810 94469 816 94521
rect 156 94349 816 94469
rect 156 94297 162 94349
rect 810 94297 816 94349
rect 156 94177 816 94297
rect 156 94125 162 94177
rect 810 94125 816 94177
rect 156 94005 816 94125
rect 156 93953 162 94005
rect 810 93953 816 94005
rect 156 93833 816 93953
rect 156 93781 162 93833
rect 810 93781 816 93833
rect 156 93661 816 93781
rect 156 93609 162 93661
rect 810 93609 816 93661
rect 156 93489 816 93609
rect 156 93437 162 93489
rect 810 93437 816 93489
rect 156 93317 816 93437
rect 156 93265 162 93317
rect 810 93265 816 93317
rect 156 93145 816 93265
rect 156 93093 162 93145
rect 810 93093 816 93145
rect 156 92973 816 93093
rect 156 92921 162 92973
rect 810 92921 816 92973
rect 156 92801 816 92921
rect 156 92749 162 92801
rect 810 92749 816 92801
rect 156 92629 816 92749
rect 156 92577 162 92629
rect 810 92577 816 92629
rect 156 92457 816 92577
rect 156 92405 162 92457
rect 810 92405 816 92457
rect 156 92285 816 92405
rect 156 92233 162 92285
rect 810 92233 816 92285
rect 156 92113 816 92233
rect 156 92061 162 92113
rect 810 92061 816 92113
rect 156 91941 816 92061
rect 156 91889 162 91941
rect 810 91889 816 91941
rect 156 91769 816 91889
rect 156 91717 162 91769
rect 810 91717 816 91769
rect 156 91597 816 91717
rect 156 91545 162 91597
rect 810 91545 816 91597
rect 156 91425 816 91545
rect 156 91373 162 91425
rect 810 91373 816 91425
rect 156 91253 816 91373
rect 156 91201 162 91253
rect 810 91201 816 91253
rect 156 91081 816 91201
rect 156 91029 162 91081
rect 810 91029 816 91081
rect 156 90909 816 91029
rect 156 90857 162 90909
rect 810 90857 816 90909
rect 156 90737 816 90857
rect 156 90685 162 90737
rect 810 90685 816 90737
rect 156 90565 816 90685
rect 156 90513 162 90565
rect 810 90513 816 90565
rect 156 90393 816 90513
rect 156 90341 162 90393
rect 810 90341 816 90393
rect 156 90221 816 90341
rect 156 90169 162 90221
rect 810 90169 816 90221
rect 156 90049 816 90169
rect 156 89997 162 90049
rect 810 89997 816 90049
rect 156 89877 816 89997
rect 156 89825 162 89877
rect 810 89825 816 89877
rect 156 89705 816 89825
rect 156 89653 162 89705
rect 810 89653 816 89705
rect 156 89533 816 89653
rect 156 89481 162 89533
rect 810 89481 816 89533
rect 156 89361 816 89481
rect 156 89309 162 89361
rect 810 89309 816 89361
rect 156 89189 816 89309
rect 156 89137 162 89189
rect 810 89137 816 89189
rect 156 89017 816 89137
rect 156 88965 162 89017
rect 810 88965 816 89017
rect 156 88845 816 88965
rect 156 88793 162 88845
rect 810 88793 816 88845
rect 156 88673 816 88793
rect 156 88621 162 88673
rect 810 88621 816 88673
rect 156 88501 816 88621
rect 156 88449 162 88501
rect 810 88449 816 88501
rect 156 88329 816 88449
rect 156 88277 162 88329
rect 810 88277 816 88329
rect 156 88157 816 88277
rect 156 88105 162 88157
rect 810 88105 816 88157
rect 156 87985 816 88105
rect 156 87933 162 87985
rect 810 87933 816 87985
rect 156 87813 816 87933
rect 156 87761 162 87813
rect 810 87761 816 87813
rect 156 87641 816 87761
rect 156 87589 162 87641
rect 810 87589 816 87641
rect 156 87469 816 87589
rect 156 87417 162 87469
rect 810 87417 816 87469
rect 156 87297 816 87417
rect 156 87245 162 87297
rect 810 87245 816 87297
rect 156 87125 816 87245
rect 156 87073 162 87125
rect 810 87073 816 87125
rect 156 86953 816 87073
rect 156 86901 162 86953
rect 810 86901 816 86953
rect 156 86781 816 86901
rect 156 86729 162 86781
rect 810 86729 816 86781
rect 156 86609 816 86729
rect 156 86557 162 86609
rect 810 86557 816 86609
rect 156 86437 816 86557
rect 156 86385 162 86437
rect 810 86385 816 86437
rect 156 86265 816 86385
rect 156 86213 162 86265
rect 810 86213 816 86265
rect 156 86093 816 86213
rect 156 86041 162 86093
rect 810 86041 816 86093
rect 156 85921 816 86041
rect 156 85869 162 85921
rect 810 85869 816 85921
rect 156 85749 816 85869
rect 156 85697 162 85749
rect 810 85697 816 85749
rect 156 85577 816 85697
rect 156 85525 162 85577
rect 810 85525 816 85577
rect 156 85405 816 85525
rect 156 85353 162 85405
rect 810 85353 816 85405
rect 156 85233 816 85353
rect 156 85181 162 85233
rect 810 85181 816 85233
rect 156 85061 816 85181
rect 156 85009 162 85061
rect 810 85009 816 85061
rect 156 84889 816 85009
rect 156 84837 162 84889
rect 810 84837 816 84889
rect 156 84717 816 84837
rect 156 84665 162 84717
rect 810 84665 816 84717
rect 156 84545 816 84665
rect 156 84493 162 84545
rect 810 84493 816 84545
rect 156 84373 816 84493
rect 156 84321 162 84373
rect 810 84321 816 84373
rect 156 84201 816 84321
rect 156 84149 162 84201
rect 810 84149 816 84201
rect 156 84029 816 84149
rect 156 83977 162 84029
rect 810 83977 816 84029
rect 156 83857 816 83977
rect 156 83805 162 83857
rect 810 83805 816 83857
rect 156 83685 816 83805
rect 156 83633 162 83685
rect 810 83633 816 83685
rect 156 83513 816 83633
rect 156 83461 162 83513
rect 810 83461 816 83513
rect 156 83341 816 83461
rect 156 83289 162 83341
rect 810 83289 816 83341
rect 156 83169 816 83289
rect 156 83117 162 83169
rect 810 83117 816 83169
rect 156 82997 816 83117
rect 156 82945 162 82997
rect 810 82945 816 82997
rect 156 82825 816 82945
rect 156 82773 162 82825
rect 810 82773 816 82825
rect 156 82653 816 82773
rect 156 82601 162 82653
rect 810 82601 816 82653
rect 156 82481 816 82601
rect 156 82429 162 82481
rect 810 82429 816 82481
rect 156 82309 816 82429
rect 156 82257 162 82309
rect 810 82257 816 82309
rect 156 82137 816 82257
rect 156 82085 162 82137
rect 810 82085 816 82137
rect 156 81965 816 82085
rect 156 81913 162 81965
rect 810 81913 816 81965
rect 156 81793 816 81913
rect 156 81741 162 81793
rect 810 81741 816 81793
rect 156 81621 816 81741
rect 156 81569 162 81621
rect 810 81569 816 81621
rect 156 81449 816 81569
rect 156 81397 162 81449
rect 810 81397 816 81449
rect 156 81277 816 81397
rect 156 81225 162 81277
rect 810 81225 816 81277
rect 156 81105 816 81225
rect 156 81053 162 81105
rect 810 81053 816 81105
rect 156 80933 816 81053
rect 156 80881 162 80933
rect 810 80881 816 80933
rect 156 80761 816 80881
rect 156 80709 162 80761
rect 810 80709 816 80761
rect 156 80589 816 80709
rect 156 80537 162 80589
rect 810 80537 816 80589
rect 156 80417 816 80537
rect 156 80365 162 80417
rect 810 80365 816 80417
rect 156 80245 816 80365
rect 156 80193 162 80245
rect 810 80193 816 80245
rect 156 80073 816 80193
rect 156 80021 162 80073
rect 810 80021 816 80073
rect 156 79901 816 80021
rect 156 79849 162 79901
rect 810 79849 816 79901
rect 156 79729 816 79849
rect 156 79677 162 79729
rect 810 79677 816 79729
rect 156 79557 816 79677
rect 156 79505 162 79557
rect 810 79505 816 79557
rect 156 79385 816 79505
rect 156 79333 162 79385
rect 810 79333 816 79385
rect 156 79213 816 79333
rect 156 79161 162 79213
rect 810 79161 816 79213
rect 156 79041 816 79161
rect 156 78989 162 79041
rect 810 78989 816 79041
rect 156 78869 816 78989
rect 156 78817 162 78869
rect 810 78817 816 78869
rect 156 78697 816 78817
rect 156 78645 162 78697
rect 810 78645 816 78697
rect 156 78525 816 78645
rect 156 78473 162 78525
rect 810 78473 816 78525
rect 156 78353 816 78473
rect 156 78301 162 78353
rect 810 78301 816 78353
rect 156 78181 816 78301
rect 156 78129 162 78181
rect 810 78129 816 78181
rect 156 78009 816 78129
rect 156 77957 162 78009
rect 810 77957 816 78009
rect 156 77837 816 77957
rect 156 77785 162 77837
rect 810 77785 816 77837
rect 156 77665 816 77785
rect 156 77613 162 77665
rect 810 77613 816 77665
rect 156 77493 816 77613
rect 156 77441 162 77493
rect 810 77441 816 77493
rect 156 77321 816 77441
rect 156 77269 162 77321
rect 810 77269 816 77321
rect 156 77149 816 77269
rect 156 77097 162 77149
rect 810 77097 816 77149
rect 156 76977 816 77097
rect 156 76925 162 76977
rect 810 76925 816 76977
rect 156 76805 816 76925
rect 156 76753 162 76805
rect 810 76753 816 76805
rect 156 76633 816 76753
rect 156 76581 162 76633
rect 810 76581 816 76633
rect 156 76461 816 76581
rect 156 76409 162 76461
rect 810 76409 816 76461
rect 156 76289 816 76409
rect 156 76237 162 76289
rect 810 76237 816 76289
rect 156 76117 816 76237
rect 156 76065 162 76117
rect 810 76065 816 76117
rect 156 75945 816 76065
rect 156 75893 162 75945
rect 810 75893 816 75945
rect 156 75773 816 75893
rect 156 75721 162 75773
rect 810 75721 816 75773
rect 156 75601 816 75721
rect 156 75549 162 75601
rect 810 75549 816 75601
rect 156 75429 816 75549
rect 156 75377 162 75429
rect 810 75377 816 75429
rect 156 75257 816 75377
rect 156 75205 162 75257
rect 810 75205 816 75257
rect 156 75085 816 75205
rect 156 75033 162 75085
rect 810 75033 816 75085
rect 156 74913 816 75033
rect 156 74861 162 74913
rect 810 74861 816 74913
rect 156 74741 816 74861
rect 156 74689 162 74741
rect 810 74689 816 74741
rect 156 74569 816 74689
rect 156 74517 162 74569
rect 810 74517 816 74569
rect 156 74397 816 74517
rect 156 74345 162 74397
rect 810 74345 816 74397
rect 156 74225 816 74345
rect 156 74173 162 74225
rect 810 74173 816 74225
rect 156 74053 816 74173
rect 156 74001 162 74053
rect 810 74001 816 74053
rect 156 73881 816 74001
rect 156 73829 162 73881
rect 810 73829 816 73881
rect 156 73709 816 73829
rect 156 73657 162 73709
rect 810 73657 816 73709
rect 156 73537 816 73657
rect 156 73485 162 73537
rect 810 73485 816 73537
rect 156 73365 816 73485
rect 156 73313 162 73365
rect 810 73313 816 73365
rect 156 73193 816 73313
rect 156 73141 162 73193
rect 810 73141 816 73193
rect 156 73021 816 73141
rect 156 72969 162 73021
rect 810 72969 816 73021
rect 156 72849 816 72969
rect 156 72797 162 72849
rect 810 72797 816 72849
rect 156 72677 816 72797
rect 156 72625 162 72677
rect 810 72625 816 72677
rect 156 72505 816 72625
rect 156 72453 162 72505
rect 810 72453 816 72505
rect 156 72333 816 72453
rect 156 72281 162 72333
rect 810 72281 816 72333
rect 156 72161 816 72281
rect 156 72109 162 72161
rect 810 72109 816 72161
rect 156 71989 816 72109
rect 156 71937 162 71989
rect 810 71937 816 71989
rect 156 71817 816 71937
rect 156 71765 162 71817
rect 810 71765 816 71817
rect 156 71645 816 71765
rect 156 71593 162 71645
rect 810 71593 816 71645
rect 156 71473 816 71593
rect 156 71421 162 71473
rect 810 71421 816 71473
rect 156 71301 816 71421
rect 156 71249 162 71301
rect 810 71249 816 71301
rect 156 71129 816 71249
rect 156 71077 162 71129
rect 810 71077 816 71129
rect 156 70957 816 71077
rect 156 70905 162 70957
rect 810 70905 816 70957
rect 156 70785 816 70905
rect 156 70733 162 70785
rect 810 70733 816 70785
rect 156 70613 816 70733
rect 156 70561 162 70613
rect 810 70561 816 70613
rect 156 70441 816 70561
rect 156 70389 162 70441
rect 810 70389 816 70441
rect 156 70269 816 70389
rect 156 70217 162 70269
rect 810 70217 816 70269
rect 156 70097 816 70217
rect 156 70045 162 70097
rect 810 70045 816 70097
rect 156 69925 816 70045
rect 156 69873 162 69925
rect 810 69873 816 69925
rect 156 69753 816 69873
rect 156 69701 162 69753
rect 810 69701 816 69753
rect 156 69581 816 69701
rect 156 69529 162 69581
rect 810 69529 816 69581
rect 156 69409 816 69529
rect 156 69357 162 69409
rect 810 69357 816 69409
rect 156 69237 816 69357
rect 156 69185 162 69237
rect 810 69185 816 69237
rect 156 69065 816 69185
rect 156 69013 162 69065
rect 810 69013 816 69065
rect 156 68893 816 69013
rect 156 68841 162 68893
rect 810 68841 816 68893
rect 156 68721 816 68841
rect 156 68669 162 68721
rect 810 68669 816 68721
rect 156 68549 816 68669
rect 156 68497 162 68549
rect 810 68497 816 68549
rect 156 68377 816 68497
rect 156 68325 162 68377
rect 810 68325 816 68377
rect 156 68205 816 68325
rect 156 68153 162 68205
rect 810 68153 816 68205
rect 156 68033 816 68153
rect 156 67981 162 68033
rect 810 67981 816 68033
rect 156 67861 816 67981
rect 156 67809 162 67861
rect 810 67809 816 67861
rect 156 67689 816 67809
rect 156 67637 162 67689
rect 810 67637 816 67689
rect 156 67517 816 67637
rect 156 67465 162 67517
rect 810 67465 816 67517
rect 156 67345 816 67465
rect 156 67293 162 67345
rect 810 67293 816 67345
rect 156 67173 816 67293
rect 156 67121 162 67173
rect 810 67121 816 67173
rect 156 67001 816 67121
rect 156 66949 162 67001
rect 810 66949 816 67001
rect 156 66829 816 66949
rect 156 66777 162 66829
rect 810 66777 816 66829
rect 156 66657 816 66777
rect 156 66605 162 66657
rect 810 66605 816 66657
rect 156 66485 816 66605
rect 156 66433 162 66485
rect 810 66433 816 66485
rect 156 66313 816 66433
rect 156 66261 162 66313
rect 810 66261 816 66313
rect 156 66141 816 66261
rect 156 66089 162 66141
rect 810 66089 816 66141
rect 156 65969 816 66089
rect 156 65917 162 65969
rect 810 65917 816 65969
rect 156 65797 816 65917
rect 156 65745 162 65797
rect 810 65745 816 65797
rect 156 65625 816 65745
rect 156 65573 162 65625
rect 810 65573 816 65625
rect 156 65453 816 65573
rect 156 65401 162 65453
rect 810 65401 816 65453
rect 156 65281 816 65401
rect 156 65229 162 65281
rect 810 65229 816 65281
rect 156 65109 816 65229
rect 156 65057 162 65109
rect 810 65057 816 65109
rect 156 64937 816 65057
rect 156 64885 162 64937
rect 810 64885 816 64937
rect 156 64765 816 64885
rect 156 64713 162 64765
rect 810 64713 816 64765
rect 156 64593 816 64713
rect 156 64541 162 64593
rect 810 64541 816 64593
rect 156 64421 816 64541
rect 156 64369 162 64421
rect 810 64369 816 64421
rect 156 64249 816 64369
rect 156 64197 162 64249
rect 810 64197 816 64249
rect 156 64077 816 64197
rect 156 64025 162 64077
rect 810 64025 816 64077
rect 156 63905 816 64025
rect 156 63853 162 63905
rect 810 63853 816 63905
rect 156 63733 816 63853
rect 156 63681 162 63733
rect 810 63681 816 63733
rect 156 63561 816 63681
rect 156 63509 162 63561
rect 810 63509 816 63561
rect 156 63389 816 63509
rect 156 63337 162 63389
rect 810 63337 816 63389
rect 156 63217 816 63337
rect 156 63165 162 63217
rect 810 63165 816 63217
rect 156 63045 816 63165
rect 156 62993 162 63045
rect 810 62993 816 63045
rect 156 62873 816 62993
rect 156 62821 162 62873
rect 810 62821 816 62873
rect 156 62701 816 62821
rect 156 62649 162 62701
rect 810 62649 816 62701
rect 156 62529 816 62649
rect 156 62477 162 62529
rect 810 62477 816 62529
rect 156 62357 816 62477
rect 156 62305 162 62357
rect 810 62305 816 62357
rect 156 62185 816 62305
rect 156 62133 162 62185
rect 810 62133 816 62185
rect 156 62013 816 62133
rect 156 61961 162 62013
rect 810 61961 816 62013
rect 156 61841 816 61961
rect 156 61789 162 61841
rect 810 61789 816 61841
rect 156 61669 816 61789
rect 156 61617 162 61669
rect 810 61617 816 61669
rect 156 61497 816 61617
rect 156 61445 162 61497
rect 810 61445 816 61497
rect 156 61325 816 61445
rect 156 61273 162 61325
rect 810 61273 816 61325
rect 156 61153 816 61273
rect 156 61101 162 61153
rect 810 61101 816 61153
rect 156 60981 816 61101
rect 156 60929 162 60981
rect 810 60929 816 60981
rect 156 60809 816 60929
rect 156 60757 162 60809
rect 810 60757 816 60809
rect 156 60637 816 60757
rect 156 60585 162 60637
rect 810 60585 816 60637
rect 156 60465 816 60585
rect 156 60413 162 60465
rect 810 60413 816 60465
rect 156 60293 816 60413
rect 156 60241 162 60293
rect 810 60241 816 60293
rect 156 60121 816 60241
rect 156 60069 162 60121
rect 810 60069 816 60121
rect 156 59949 816 60069
rect 156 59897 162 59949
rect 810 59897 816 59949
rect 156 59777 816 59897
rect 156 59725 162 59777
rect 810 59725 816 59777
rect 156 59605 816 59725
rect 156 59553 162 59605
rect 810 59553 816 59605
rect 156 59433 816 59553
rect 156 59381 162 59433
rect 810 59381 816 59433
rect 156 59261 816 59381
rect 156 59209 162 59261
rect 810 59209 816 59261
rect 156 59089 816 59209
rect 156 59037 162 59089
rect 810 59037 816 59089
rect 156 58917 816 59037
rect 156 58865 162 58917
rect 810 58865 816 58917
rect 156 58745 816 58865
rect 156 58693 162 58745
rect 810 58693 816 58745
rect 156 58573 816 58693
rect 156 58521 162 58573
rect 810 58521 816 58573
rect 156 58401 816 58521
rect 156 58349 162 58401
rect 810 58349 816 58401
rect 156 58229 816 58349
rect 156 58177 162 58229
rect 810 58177 816 58229
rect 156 58057 816 58177
rect 156 58005 162 58057
rect 810 58005 816 58057
rect 156 57885 816 58005
rect 156 57833 162 57885
rect 810 57833 816 57885
rect 156 57713 816 57833
rect 156 57661 162 57713
rect 810 57661 816 57713
rect 156 57541 816 57661
rect 156 57489 162 57541
rect 810 57489 816 57541
rect 156 57369 816 57489
rect 156 57317 162 57369
rect 810 57317 816 57369
rect 156 57197 816 57317
rect 156 57145 162 57197
rect 810 57145 816 57197
rect 156 57025 816 57145
rect 156 56973 162 57025
rect 810 56973 816 57025
rect 156 56853 816 56973
rect 156 56801 162 56853
rect 810 56801 816 56853
rect 156 56681 816 56801
rect 156 56629 162 56681
rect 810 56629 816 56681
rect 156 56509 816 56629
rect 156 56457 162 56509
rect 810 56457 816 56509
rect 156 56337 816 56457
rect 156 56285 162 56337
rect 810 56285 816 56337
rect 156 56165 816 56285
rect 156 56113 162 56165
rect 810 56113 816 56165
rect 156 55993 816 56113
rect 156 55941 162 55993
rect 810 55941 816 55993
rect 156 55821 816 55941
rect 156 55769 162 55821
rect 810 55769 816 55821
rect 156 55649 816 55769
rect 156 55597 162 55649
rect 810 55597 816 55649
rect 156 55477 816 55597
rect 156 55425 162 55477
rect 810 55425 816 55477
rect 156 55305 816 55425
rect 156 55253 162 55305
rect 810 55253 816 55305
rect 156 55133 816 55253
rect 156 55081 162 55133
rect 810 55081 816 55133
rect 156 54961 816 55081
rect 156 54909 162 54961
rect 810 54909 816 54961
rect 156 54789 816 54909
rect 156 54737 162 54789
rect 810 54737 816 54789
rect 156 54617 816 54737
rect 156 54565 162 54617
rect 810 54565 816 54617
rect 156 54445 816 54565
rect 156 54393 162 54445
rect 810 54393 816 54445
rect 156 54273 816 54393
rect 156 54221 162 54273
rect 810 54221 816 54273
rect 156 54101 816 54221
rect 156 54049 162 54101
rect 810 54049 816 54101
rect 156 53929 816 54049
rect 156 53877 162 53929
rect 810 53877 816 53929
rect 156 53757 816 53877
rect 156 53705 162 53757
rect 810 53705 816 53757
rect 156 53585 816 53705
rect 156 53533 162 53585
rect 810 53533 816 53585
rect 156 53413 816 53533
rect 156 53361 162 53413
rect 810 53361 816 53413
rect 156 53241 816 53361
rect 156 53189 162 53241
rect 810 53189 816 53241
rect 156 53069 816 53189
rect 156 53017 162 53069
rect 810 53017 816 53069
rect 156 52897 816 53017
rect 156 52845 162 52897
rect 810 52845 816 52897
rect 156 52725 816 52845
rect 156 52673 162 52725
rect 810 52673 816 52725
rect 156 52553 816 52673
rect 156 52501 162 52553
rect 810 52501 816 52553
rect 156 52381 816 52501
rect 156 52329 162 52381
rect 810 52329 816 52381
rect 156 52209 816 52329
rect 156 52157 162 52209
rect 810 52157 816 52209
rect 156 52037 816 52157
rect 156 51985 162 52037
rect 810 51985 816 52037
rect 156 51865 816 51985
rect 156 51813 162 51865
rect 810 51813 816 51865
rect 156 51693 816 51813
rect 156 51641 162 51693
rect 810 51641 816 51693
rect 156 51521 816 51641
rect 156 51469 162 51521
rect 810 51469 816 51521
rect 156 51349 816 51469
rect 156 51297 162 51349
rect 810 51297 816 51349
rect 156 51177 816 51297
rect 156 51125 162 51177
rect 810 51125 816 51177
rect 156 51005 816 51125
rect 156 50953 162 51005
rect 810 50953 816 51005
rect 156 50833 816 50953
rect 156 50781 162 50833
rect 810 50781 816 50833
rect 156 50661 816 50781
rect 156 50609 162 50661
rect 810 50609 816 50661
rect 156 50489 816 50609
rect 156 50437 162 50489
rect 810 50437 816 50489
rect 156 50317 816 50437
rect 156 50265 162 50317
rect 810 50265 816 50317
rect 156 50145 816 50265
rect 156 50093 162 50145
rect 810 50093 816 50145
rect 156 49973 816 50093
rect 156 49921 162 49973
rect 810 49921 816 49973
rect 156 49801 816 49921
rect 156 49749 162 49801
rect 810 49749 816 49801
rect 156 49629 816 49749
rect 156 49577 162 49629
rect 810 49577 816 49629
rect 156 49457 816 49577
rect 156 49405 162 49457
rect 810 49405 816 49457
rect 156 49285 816 49405
rect 156 49233 162 49285
rect 810 49233 816 49285
rect 156 49113 816 49233
rect 156 49061 162 49113
rect 810 49061 816 49113
rect 156 48941 816 49061
rect 156 48889 162 48941
rect 810 48889 816 48941
rect 156 48769 816 48889
rect 156 48717 162 48769
rect 810 48717 816 48769
rect 156 48597 816 48717
rect 156 48545 162 48597
rect 810 48545 816 48597
rect 156 48425 816 48545
rect 156 48373 162 48425
rect 810 48373 816 48425
rect 156 48253 816 48373
rect 156 48201 162 48253
rect 810 48201 816 48253
rect 156 48081 816 48201
rect 156 48029 162 48081
rect 810 48029 816 48081
rect 156 47909 816 48029
rect 156 47857 162 47909
rect 810 47857 816 47909
rect 156 47737 816 47857
rect 156 47685 162 47737
rect 810 47685 816 47737
rect 156 47565 816 47685
rect 156 47513 162 47565
rect 810 47513 816 47565
rect 156 47393 816 47513
rect 156 47341 162 47393
rect 810 47341 816 47393
rect 156 47221 816 47341
rect 156 47169 162 47221
rect 810 47169 816 47221
rect 156 47049 816 47169
rect 156 46997 162 47049
rect 810 46997 816 47049
rect 156 46877 816 46997
rect 156 46825 162 46877
rect 810 46825 816 46877
rect 156 46705 816 46825
rect 156 46653 162 46705
rect 810 46653 816 46705
rect 156 46533 816 46653
rect 156 46481 162 46533
rect 810 46481 816 46533
rect 156 46361 816 46481
rect 156 46309 162 46361
rect 810 46309 816 46361
rect 156 46189 816 46309
rect 156 46137 162 46189
rect 810 46137 816 46189
rect 156 46017 816 46137
rect 156 45965 162 46017
rect 810 45965 816 46017
rect 156 45845 816 45965
rect 156 45793 162 45845
rect 810 45793 816 45845
rect 156 45673 816 45793
rect 156 45621 162 45673
rect 810 45621 816 45673
rect 156 45501 816 45621
rect 156 45449 162 45501
rect 810 45449 816 45501
rect 156 45329 816 45449
rect 156 45277 162 45329
rect 810 45277 816 45329
rect 156 45157 816 45277
rect 156 45105 162 45157
rect 810 45105 816 45157
rect 156 44985 816 45105
rect 156 44933 162 44985
rect 810 44933 816 44985
rect 156 44813 816 44933
rect 156 44761 162 44813
rect 810 44761 816 44813
rect 156 44641 816 44761
rect 156 44589 162 44641
rect 810 44589 816 44641
rect 156 44469 816 44589
rect 156 44417 162 44469
rect 810 44417 816 44469
rect 156 44297 816 44417
rect 156 44245 162 44297
rect 810 44245 816 44297
rect 156 44125 816 44245
rect 156 44073 162 44125
rect 810 44073 816 44125
rect 156 43953 816 44073
rect 156 43901 162 43953
rect 810 43901 816 43953
rect 156 43781 816 43901
rect 156 43729 162 43781
rect 810 43729 816 43781
rect 156 43609 816 43729
rect 156 43557 162 43609
rect 810 43557 816 43609
rect 156 43437 816 43557
rect 156 43385 162 43437
rect 810 43385 816 43437
rect 156 43265 816 43385
rect 156 43213 162 43265
rect 810 43213 816 43265
rect 156 43093 816 43213
rect 156 43041 162 43093
rect 810 43041 816 43093
rect 156 42921 816 43041
rect 156 42869 162 42921
rect 810 42869 816 42921
rect 156 42749 816 42869
rect 156 42697 162 42749
rect 810 42697 816 42749
rect 156 42577 816 42697
rect 156 42525 162 42577
rect 810 42525 816 42577
rect 156 42405 816 42525
rect 156 42353 162 42405
rect 810 42353 816 42405
rect 156 42233 816 42353
rect 156 42181 162 42233
rect 810 42181 816 42233
rect 156 42061 816 42181
rect 156 42009 162 42061
rect 810 42009 816 42061
rect 156 41889 816 42009
rect 156 41837 162 41889
rect 810 41837 816 41889
rect 156 41717 816 41837
rect 156 41665 162 41717
rect 810 41665 816 41717
rect 156 41545 816 41665
rect 156 41493 162 41545
rect 810 41493 816 41545
rect 156 41373 816 41493
rect 156 41321 162 41373
rect 810 41321 816 41373
rect 156 41201 816 41321
rect 156 41149 162 41201
rect 810 41149 816 41201
rect 156 41029 816 41149
rect 156 40977 162 41029
rect 810 40977 816 41029
rect 156 40857 816 40977
rect 156 40805 162 40857
rect 810 40805 816 40857
rect 156 40685 816 40805
rect 156 40633 162 40685
rect 810 40633 816 40685
rect 156 40513 816 40633
rect 156 40461 162 40513
rect 810 40461 816 40513
rect 156 40341 816 40461
rect 156 40289 162 40341
rect 810 40289 816 40341
rect 156 40169 816 40289
rect 156 40117 162 40169
rect 810 40117 816 40169
rect 156 39997 816 40117
rect 156 39945 162 39997
rect 810 39945 816 39997
rect 156 39825 816 39945
rect 156 39773 162 39825
rect 810 39773 816 39825
rect 156 39653 816 39773
rect 156 39601 162 39653
rect 810 39601 816 39653
rect 156 39481 816 39601
rect 156 39429 162 39481
rect 810 39429 816 39481
rect 156 39309 816 39429
rect 156 39257 162 39309
rect 810 39257 816 39309
rect 156 39137 816 39257
rect 156 39085 162 39137
rect 810 39085 816 39137
rect 156 38965 816 39085
rect 156 38913 162 38965
rect 810 38913 816 38965
rect 156 38793 816 38913
rect 156 38741 162 38793
rect 810 38741 816 38793
rect 156 38621 816 38741
rect 156 38569 162 38621
rect 810 38569 816 38621
rect 156 38449 816 38569
rect 156 38397 162 38449
rect 810 38397 816 38449
rect 156 38277 816 38397
rect 156 38225 162 38277
rect 810 38225 816 38277
rect 156 38105 816 38225
rect 156 38053 162 38105
rect 810 38053 816 38105
rect 156 37933 816 38053
rect 156 37881 162 37933
rect 810 37881 816 37933
rect 156 37761 816 37881
rect 156 37709 162 37761
rect 810 37709 816 37761
rect 156 37589 816 37709
rect 156 37537 162 37589
rect 810 37537 816 37589
rect 156 37417 816 37537
rect 156 37365 162 37417
rect 810 37365 816 37417
rect 156 37245 816 37365
rect 156 37193 162 37245
rect 810 37193 816 37245
rect 156 37073 816 37193
rect 156 37021 162 37073
rect 810 37021 816 37073
rect 156 36901 816 37021
rect 156 36849 162 36901
rect 810 36849 816 36901
rect 156 36729 816 36849
rect 156 36677 162 36729
rect 810 36677 816 36729
rect 156 36557 816 36677
rect 156 36505 162 36557
rect 810 36505 816 36557
rect 156 36385 816 36505
rect 156 36333 162 36385
rect 810 36333 816 36385
rect 156 36213 816 36333
rect 156 36161 162 36213
rect 810 36161 816 36213
rect 156 36041 816 36161
rect 156 35989 162 36041
rect 810 35989 816 36041
rect 156 35869 816 35989
rect 156 35817 162 35869
rect 810 35817 816 35869
rect 156 35697 816 35817
rect 156 35645 162 35697
rect 810 35645 816 35697
rect 156 35525 816 35645
rect 156 35473 162 35525
rect 810 35473 816 35525
rect 156 35353 816 35473
rect 156 35301 162 35353
rect 810 35301 816 35353
rect 156 35181 816 35301
rect 156 35129 162 35181
rect 810 35129 816 35181
rect 156 35009 816 35129
rect 156 34957 162 35009
rect 810 34957 816 35009
rect 156 34837 816 34957
rect 156 34785 162 34837
rect 810 34785 816 34837
rect 156 34665 816 34785
rect 156 34613 162 34665
rect 810 34613 816 34665
rect 156 34493 816 34613
rect 156 34441 162 34493
rect 810 34441 816 34493
rect 156 34321 816 34441
rect 156 34269 162 34321
rect 810 34269 816 34321
rect 156 34149 816 34269
rect 156 34097 162 34149
rect 810 34097 816 34149
rect 156 33977 816 34097
rect 156 33925 162 33977
rect 810 33925 816 33977
rect 156 33805 816 33925
rect 156 33753 162 33805
rect 810 33753 816 33805
rect 156 33633 816 33753
rect 156 33581 162 33633
rect 810 33581 816 33633
rect 156 33461 816 33581
rect 156 33409 162 33461
rect 810 33409 816 33461
rect 156 33289 816 33409
rect 156 33237 162 33289
rect 810 33237 816 33289
rect 156 33117 816 33237
rect 156 33065 162 33117
rect 810 33065 816 33117
rect 156 32945 816 33065
rect 156 32893 162 32945
rect 810 32893 816 32945
rect 156 32773 816 32893
rect 156 32721 162 32773
rect 810 32721 816 32773
rect 156 32601 816 32721
rect 156 32549 162 32601
rect 810 32549 816 32601
rect 156 32429 816 32549
rect 156 32377 162 32429
rect 810 32377 816 32429
rect 156 32257 816 32377
rect 156 32205 162 32257
rect 810 32205 816 32257
rect 156 32085 816 32205
rect 156 32033 162 32085
rect 810 32033 816 32085
rect 156 31913 816 32033
rect 156 31861 162 31913
rect 810 31861 816 31913
rect 156 31741 816 31861
rect 156 31689 162 31741
rect 810 31689 816 31741
rect 156 31569 816 31689
rect 156 31517 162 31569
rect 810 31517 816 31569
rect 156 31397 816 31517
rect 156 31345 162 31397
rect 810 31345 816 31397
rect 156 31225 816 31345
rect 156 31173 162 31225
rect 810 31173 816 31225
rect 156 31053 816 31173
rect 156 31001 162 31053
rect 810 31001 816 31053
rect 156 30881 816 31001
rect 156 30829 162 30881
rect 810 30829 816 30881
rect 156 30709 816 30829
rect 156 30657 162 30709
rect 810 30657 816 30709
rect 156 30537 816 30657
rect 156 30485 162 30537
rect 810 30485 816 30537
rect 156 30365 816 30485
rect 156 30313 162 30365
rect 810 30313 816 30365
rect 156 30193 816 30313
rect 156 30141 162 30193
rect 810 30141 816 30193
rect 156 30021 816 30141
rect 156 29969 162 30021
rect 810 29969 816 30021
rect 156 29849 816 29969
rect 156 29797 162 29849
rect 810 29797 816 29849
rect 156 29677 816 29797
rect 156 29625 162 29677
rect 810 29625 816 29677
rect 156 29505 816 29625
rect 156 29453 162 29505
rect 810 29453 816 29505
rect 156 29333 816 29453
rect 156 29281 162 29333
rect 810 29281 816 29333
rect 156 29161 816 29281
rect 156 29109 162 29161
rect 810 29109 816 29161
rect 156 28989 816 29109
rect 156 28937 162 28989
rect 810 28937 816 28989
rect 156 28817 816 28937
rect 156 28765 162 28817
rect 810 28765 816 28817
rect 156 28645 816 28765
rect 156 28593 162 28645
rect 810 28593 816 28645
rect 156 28473 816 28593
rect 156 28421 162 28473
rect 810 28421 816 28473
rect 156 28301 816 28421
rect 156 28249 162 28301
rect 810 28249 816 28301
rect 156 28129 816 28249
rect 156 28077 162 28129
rect 810 28077 816 28129
rect 156 27957 816 28077
rect 156 27905 162 27957
rect 810 27905 816 27957
rect 156 27785 816 27905
rect 156 27733 162 27785
rect 810 27733 816 27785
rect 156 27613 816 27733
rect 156 27561 162 27613
rect 810 27561 816 27613
rect 156 27441 816 27561
rect 156 27389 162 27441
rect 810 27389 816 27441
rect 156 27269 816 27389
rect 156 27217 162 27269
rect 810 27217 816 27269
rect 156 27097 816 27217
rect 156 27045 162 27097
rect 810 27045 816 27097
rect 156 26925 816 27045
rect 156 26873 162 26925
rect 810 26873 816 26925
rect 156 26753 816 26873
rect 156 26701 162 26753
rect 810 26701 816 26753
rect 156 26581 816 26701
rect 156 26529 162 26581
rect 810 26529 816 26581
rect 156 26409 816 26529
rect 156 26357 162 26409
rect 810 26357 816 26409
rect 156 26237 816 26357
rect 156 26185 162 26237
rect 810 26185 816 26237
rect 156 26065 816 26185
rect 156 26013 162 26065
rect 810 26013 816 26065
rect 156 25893 816 26013
rect 156 25841 162 25893
rect 810 25841 816 25893
rect 156 25721 816 25841
rect 156 25669 162 25721
rect 810 25669 816 25721
rect 156 25549 816 25669
rect 156 25497 162 25549
rect 810 25497 816 25549
rect 156 25377 816 25497
rect 156 25325 162 25377
rect 810 25325 816 25377
rect 156 25205 816 25325
rect 156 25153 162 25205
rect 810 25153 816 25205
rect 156 25033 816 25153
rect 156 24981 162 25033
rect 810 24981 816 25033
rect 156 24861 816 24981
rect 156 24809 162 24861
rect 810 24809 816 24861
rect 156 24689 816 24809
rect 156 24637 162 24689
rect 810 24637 816 24689
rect 156 24517 816 24637
rect 156 24465 162 24517
rect 810 24465 816 24517
rect 156 24345 816 24465
rect 156 24293 162 24345
rect 810 24293 816 24345
rect 156 24173 816 24293
rect 156 24121 162 24173
rect 810 24121 816 24173
rect 156 24001 816 24121
rect 156 23949 162 24001
rect 810 23949 816 24001
rect 156 23829 816 23949
rect 156 23777 162 23829
rect 810 23777 816 23829
rect 156 23657 816 23777
rect 156 23605 162 23657
rect 810 23605 816 23657
rect 156 23485 816 23605
rect 156 23433 162 23485
rect 810 23433 816 23485
rect 156 23313 816 23433
rect 156 23261 162 23313
rect 810 23261 816 23313
rect 156 23141 816 23261
rect 156 23089 162 23141
rect 810 23089 816 23141
rect 156 22969 816 23089
rect 156 22917 162 22969
rect 810 22917 816 22969
rect 156 22797 816 22917
rect 156 22745 162 22797
rect 810 22745 816 22797
rect 156 22625 816 22745
rect 156 22573 162 22625
rect 810 22573 816 22625
rect 156 22453 816 22573
rect 156 22401 162 22453
rect 810 22401 816 22453
rect 156 22281 816 22401
rect 156 22229 162 22281
rect 810 22229 816 22281
rect 156 22109 816 22229
rect 156 22057 162 22109
rect 810 22057 816 22109
rect 156 21937 816 22057
rect 156 21885 162 21937
rect 810 21885 816 21937
rect 156 21765 816 21885
rect 156 21713 162 21765
rect 810 21713 816 21765
rect 156 21593 816 21713
rect 156 21541 162 21593
rect 810 21541 816 21593
rect 156 21421 816 21541
rect 156 21369 162 21421
rect 810 21369 816 21421
rect 156 21249 816 21369
rect 156 21197 162 21249
rect 810 21197 816 21249
rect 156 21077 816 21197
rect 156 21025 162 21077
rect 810 21025 816 21077
rect 156 20905 816 21025
rect 156 20853 162 20905
rect 810 20853 816 20905
rect 156 20733 816 20853
rect 156 20681 162 20733
rect 810 20681 816 20733
rect 156 20561 816 20681
rect 156 20509 162 20561
rect 810 20509 816 20561
rect 156 20389 816 20509
rect 156 20337 162 20389
rect 810 20337 816 20389
rect 156 20217 816 20337
rect 156 20165 162 20217
rect 810 20165 816 20217
rect 156 20045 816 20165
rect 156 19993 162 20045
rect 810 19993 816 20045
rect 156 19873 816 19993
rect 156 19821 162 19873
rect 810 19821 816 19873
rect 156 19701 816 19821
rect 156 19649 162 19701
rect 810 19649 816 19701
rect 156 19529 816 19649
rect 156 19477 162 19529
rect 810 19477 816 19529
rect 156 19357 816 19477
rect 156 19305 162 19357
rect 810 19305 816 19357
rect 156 19185 816 19305
rect 156 19133 162 19185
rect 810 19133 816 19185
rect 156 19013 816 19133
rect 156 18961 162 19013
rect 810 18961 816 19013
rect 156 18841 816 18961
rect 156 18789 162 18841
rect 810 18789 816 18841
rect 156 18669 816 18789
rect 156 18617 162 18669
rect 810 18617 816 18669
rect 156 18497 816 18617
rect 156 18445 162 18497
rect 810 18445 816 18497
rect 156 18325 816 18445
rect 156 18273 162 18325
rect 810 18273 816 18325
rect 156 18153 816 18273
rect 156 18101 162 18153
rect 810 18101 816 18153
rect 156 17981 816 18101
rect 156 17929 162 17981
rect 810 17929 816 17981
rect 156 17809 816 17929
rect 156 17757 162 17809
rect 810 17757 816 17809
rect 156 17637 816 17757
rect 156 17585 162 17637
rect 810 17585 816 17637
rect 156 17465 816 17585
rect 156 17413 162 17465
rect 810 17413 816 17465
rect 156 17293 816 17413
rect 156 17241 162 17293
rect 810 17241 816 17293
rect 156 17121 816 17241
rect 156 17069 162 17121
rect 810 17069 816 17121
rect 156 16949 816 17069
rect 156 16897 162 16949
rect 810 16897 816 16949
rect 156 16777 816 16897
rect 156 16725 162 16777
rect 810 16725 816 16777
rect 156 16605 816 16725
rect 156 16553 162 16605
rect 810 16553 816 16605
rect 156 16433 816 16553
rect 156 16381 162 16433
rect 810 16381 816 16433
rect 156 16261 816 16381
rect 156 16209 162 16261
rect 810 16209 816 16261
rect 156 16089 816 16209
rect 156 16037 162 16089
rect 810 16037 816 16089
rect 156 15917 816 16037
rect 156 15865 162 15917
rect 810 15865 816 15917
rect 156 15745 816 15865
rect 156 15693 162 15745
rect 810 15693 816 15745
rect 156 15573 816 15693
rect 156 15521 162 15573
rect 810 15521 816 15573
rect 156 15401 816 15521
rect 156 15349 162 15401
rect 810 15349 816 15401
rect 156 15229 816 15349
rect 156 15177 162 15229
rect 810 15177 816 15229
rect 156 15057 816 15177
rect 156 15005 162 15057
rect 810 15005 816 15057
rect 156 14885 816 15005
rect 156 14833 162 14885
rect 810 14833 816 14885
rect 156 14713 816 14833
rect 156 14661 162 14713
rect 810 14661 816 14713
rect 156 14541 816 14661
rect 156 14489 162 14541
rect 810 14489 816 14541
rect 156 14369 816 14489
rect 156 14317 162 14369
rect 810 14317 816 14369
rect 156 14197 816 14317
rect 156 14145 162 14197
rect 810 14145 816 14197
rect 156 14025 816 14145
rect 156 13973 162 14025
rect 810 13973 816 14025
rect 156 13853 816 13973
rect 156 13801 162 13853
rect 810 13801 816 13853
rect 156 13681 816 13801
rect 156 13629 162 13681
rect 810 13629 816 13681
rect 156 13509 816 13629
rect 156 13457 162 13509
rect 810 13457 816 13509
rect 156 13337 816 13457
rect 156 13285 162 13337
rect 810 13285 816 13337
rect 156 13165 816 13285
rect 156 13113 162 13165
rect 810 13113 816 13165
rect 156 12993 816 13113
rect 156 12941 162 12993
rect 810 12941 816 12993
rect 156 12821 816 12941
rect 156 12769 162 12821
rect 810 12769 816 12821
rect 156 12649 816 12769
rect 156 12597 162 12649
rect 810 12597 816 12649
rect 156 12477 816 12597
rect 156 12425 162 12477
rect 810 12425 816 12477
rect 156 12305 816 12425
rect 156 12253 162 12305
rect 810 12253 816 12305
rect 156 12133 816 12253
rect 156 12081 162 12133
rect 810 12081 816 12133
rect 156 11961 816 12081
rect 156 11909 162 11961
rect 810 11909 816 11961
rect 156 11789 816 11909
rect 156 11737 162 11789
rect 810 11737 816 11789
rect 156 11617 816 11737
rect 156 11565 162 11617
rect 810 11565 816 11617
rect 156 11445 816 11565
rect 156 11393 162 11445
rect 810 11393 816 11445
rect 156 11273 816 11393
rect 156 11221 162 11273
rect 810 11221 816 11273
rect 156 11101 816 11221
rect 156 11049 162 11101
rect 810 11049 816 11101
rect 156 10929 816 11049
rect 156 10877 162 10929
rect 810 10877 816 10929
rect 156 10757 816 10877
rect 156 10705 162 10757
rect 810 10705 816 10757
rect 156 10585 816 10705
rect 156 10533 162 10585
rect 810 10533 816 10585
rect 156 10413 816 10533
rect 156 10361 162 10413
rect 810 10361 816 10413
rect 156 10241 816 10361
rect 156 10189 162 10241
rect 810 10189 816 10241
rect 156 10069 816 10189
rect 156 10017 162 10069
rect 810 10017 816 10069
rect 156 9897 816 10017
rect 156 9845 162 9897
rect 810 9845 816 9897
rect 156 9725 816 9845
rect 156 9673 162 9725
rect 810 9673 816 9725
rect 156 9553 816 9673
rect 156 9501 162 9553
rect 810 9501 816 9553
rect 156 9381 816 9501
rect 156 9329 162 9381
rect 810 9329 816 9381
rect 156 9209 816 9329
rect 156 9157 162 9209
rect 810 9157 816 9209
rect 156 9037 816 9157
rect 156 8985 162 9037
rect 810 8985 816 9037
rect 156 8865 816 8985
rect 156 8813 162 8865
rect 810 8813 816 8865
rect 156 8693 816 8813
rect 156 8641 162 8693
rect 810 8641 816 8693
rect 156 8521 816 8641
rect 156 8469 162 8521
rect 810 8469 816 8521
rect 156 8349 816 8469
rect 156 8297 162 8349
rect 810 8297 816 8349
rect 156 8177 816 8297
rect 156 8125 162 8177
rect 810 8125 816 8177
rect 156 8005 816 8125
rect 156 7953 162 8005
rect 810 7953 816 8005
rect 156 7833 816 7953
rect 156 7781 162 7833
rect 810 7781 816 7833
rect 156 7661 816 7781
rect 156 7609 162 7661
rect 810 7609 816 7661
rect 156 7489 816 7609
rect 156 7437 162 7489
rect 810 7437 816 7489
rect 156 7317 816 7437
rect 156 7265 162 7317
rect 810 7265 816 7317
rect 156 7145 816 7265
rect 156 7093 162 7145
rect 810 7093 816 7145
rect 156 6973 816 7093
rect 156 6921 162 6973
rect 810 6921 816 6973
rect 156 6801 816 6921
rect 156 6749 162 6801
rect 810 6749 816 6801
rect 156 6629 816 6749
rect 156 6577 162 6629
rect 810 6577 816 6629
rect 156 6457 816 6577
rect 156 6405 162 6457
rect 810 6405 816 6457
rect 156 6285 816 6405
rect 156 6233 162 6285
rect 810 6233 816 6285
rect 156 6113 816 6233
rect 156 6061 162 6113
rect 810 6061 816 6113
rect 156 5941 816 6061
rect 156 5889 162 5941
rect 810 5889 816 5941
rect 156 5769 816 5889
rect 156 5717 162 5769
rect 810 5717 816 5769
rect 156 5597 816 5717
rect 156 5545 162 5597
rect 810 5545 816 5597
rect 156 5425 816 5545
rect 156 5373 162 5425
rect 810 5373 816 5425
rect 156 5253 816 5373
rect 156 5201 162 5253
rect 810 5201 816 5253
rect 156 5081 816 5201
rect 156 5029 162 5081
rect 810 5029 816 5081
rect 156 4909 816 5029
rect 156 4857 162 4909
rect 810 4857 816 4909
rect 156 4737 816 4857
rect 156 4685 162 4737
rect 810 4685 816 4737
rect 156 4565 816 4685
rect 156 4513 162 4565
rect 810 4513 816 4565
rect 156 4393 816 4513
rect 156 4341 162 4393
rect 810 4341 816 4393
rect 156 4221 816 4341
rect 156 4169 162 4221
rect 810 4169 816 4221
rect 156 4049 816 4169
rect 156 3997 162 4049
rect 810 3997 816 4049
rect 156 3877 816 3997
rect 156 3825 162 3877
rect 810 3825 816 3877
rect 156 3705 816 3825
rect 156 3653 162 3705
rect 810 3653 816 3705
rect 156 3533 816 3653
rect 156 3481 162 3533
rect 810 3481 816 3533
rect 156 3361 816 3481
rect 156 3309 162 3361
rect 810 3309 816 3361
rect 156 3189 816 3309
rect 156 3137 162 3189
rect 810 3137 816 3189
rect 156 3017 816 3137
rect 156 2965 162 3017
rect 810 2965 816 3017
rect 156 2845 816 2965
rect 156 2793 162 2845
rect 810 2793 816 2845
rect 156 2673 816 2793
rect 156 2621 162 2673
rect 810 2621 816 2673
rect 156 2501 816 2621
rect 156 2449 162 2501
rect 810 2449 816 2501
rect 156 2329 816 2449
rect 156 2277 162 2329
rect 810 2277 816 2329
rect 156 2157 816 2277
rect 156 2105 162 2157
rect 810 2105 816 2157
rect 156 1985 816 2105
rect 156 1933 162 1985
rect 810 1933 816 1985
rect 156 1813 816 1933
rect 156 1761 162 1813
rect 810 1761 816 1813
rect 156 1641 816 1761
rect 156 1589 162 1641
rect 810 1589 816 1641
rect 156 1469 816 1589
rect 156 1417 162 1469
rect 810 1417 816 1469
rect 156 1297 816 1417
rect 156 1245 162 1297
rect 810 1245 816 1297
rect 156 1125 816 1245
rect 156 1073 162 1125
rect 810 1073 816 1125
rect 156 953 816 1073
rect 156 901 162 953
rect 810 901 816 953
rect 156 781 816 901
rect 156 729 162 781
rect 810 729 816 781
rect 156 609 816 729
rect 156 557 162 609
rect 810 557 816 609
rect 156 437 816 557
rect 156 385 162 437
rect 810 385 816 437
rect 156 265 816 385
rect 156 213 162 265
rect 810 213 816 265
rect 156 127 816 213
rect 894 100059 900 100111
rect 1548 100059 1554 100111
rect 894 99939 1554 100059
rect 894 99887 900 99939
rect 1548 99887 1554 99939
rect 894 99767 1554 99887
rect 894 99715 900 99767
rect 1548 99715 1554 99767
rect 894 99595 1554 99715
rect 894 99543 900 99595
rect 1548 99543 1554 99595
rect 894 99423 1554 99543
rect 894 99371 900 99423
rect 1548 99371 1554 99423
rect 894 99251 1554 99371
rect 894 99199 900 99251
rect 1548 99199 1554 99251
rect 894 99079 1554 99199
rect 894 99027 900 99079
rect 1548 99027 1554 99079
rect 894 98907 1554 99027
rect 894 98855 900 98907
rect 1548 98855 1554 98907
rect 894 98735 1554 98855
rect 894 98683 900 98735
rect 1548 98683 1554 98735
rect 894 98563 1554 98683
rect 894 98511 900 98563
rect 1548 98511 1554 98563
rect 894 98391 1554 98511
rect 894 98339 900 98391
rect 1548 98339 1554 98391
rect 894 98219 1554 98339
rect 894 98167 900 98219
rect 1548 98167 1554 98219
rect 894 98047 1554 98167
rect 894 97995 900 98047
rect 1548 97995 1554 98047
rect 894 97875 1554 97995
rect 894 97823 900 97875
rect 1548 97823 1554 97875
rect 894 97703 1554 97823
rect 894 97651 900 97703
rect 1548 97651 1554 97703
rect 894 97531 1554 97651
rect 894 97479 900 97531
rect 1548 97479 1554 97531
rect 894 97359 1554 97479
rect 894 97307 900 97359
rect 1548 97307 1554 97359
rect 894 97187 1554 97307
rect 894 97135 900 97187
rect 1548 97135 1554 97187
rect 894 97015 1554 97135
rect 894 96963 900 97015
rect 1548 96963 1554 97015
rect 894 96843 1554 96963
rect 894 96791 900 96843
rect 1548 96791 1554 96843
rect 894 96671 1554 96791
rect 894 96619 900 96671
rect 1548 96619 1554 96671
rect 894 96499 1554 96619
rect 894 96447 900 96499
rect 1548 96447 1554 96499
rect 894 96327 1554 96447
rect 894 96275 900 96327
rect 1548 96275 1554 96327
rect 894 96155 1554 96275
rect 894 96103 900 96155
rect 1548 96103 1554 96155
rect 894 95983 1554 96103
rect 894 95931 900 95983
rect 1548 95931 1554 95983
rect 894 95811 1554 95931
rect 894 95759 900 95811
rect 1548 95759 1554 95811
rect 894 95639 1554 95759
rect 894 95587 900 95639
rect 1548 95587 1554 95639
rect 894 95467 1554 95587
rect 894 95415 900 95467
rect 1548 95415 1554 95467
rect 894 95295 1554 95415
rect 894 95243 900 95295
rect 1548 95243 1554 95295
rect 894 95123 1554 95243
rect 894 95071 900 95123
rect 1548 95071 1554 95123
rect 894 94951 1554 95071
rect 894 94899 900 94951
rect 1548 94899 1554 94951
rect 894 94779 1554 94899
rect 894 94727 900 94779
rect 1548 94727 1554 94779
rect 894 94607 1554 94727
rect 894 94555 900 94607
rect 1548 94555 1554 94607
rect 894 94435 1554 94555
rect 894 94383 900 94435
rect 1548 94383 1554 94435
rect 894 94263 1554 94383
rect 894 94211 900 94263
rect 1548 94211 1554 94263
rect 894 94091 1554 94211
rect 894 94039 900 94091
rect 1548 94039 1554 94091
rect 894 93919 1554 94039
rect 894 93867 900 93919
rect 1548 93867 1554 93919
rect 894 93747 1554 93867
rect 894 93695 900 93747
rect 1548 93695 1554 93747
rect 894 93575 1554 93695
rect 894 93523 900 93575
rect 1548 93523 1554 93575
rect 894 93403 1554 93523
rect 894 93351 900 93403
rect 1548 93351 1554 93403
rect 894 93231 1554 93351
rect 894 93179 900 93231
rect 1548 93179 1554 93231
rect 894 93059 1554 93179
rect 894 93007 900 93059
rect 1548 93007 1554 93059
rect 894 92887 1554 93007
rect 894 92835 900 92887
rect 1548 92835 1554 92887
rect 894 92715 1554 92835
rect 894 92663 900 92715
rect 1548 92663 1554 92715
rect 894 92543 1554 92663
rect 894 92491 900 92543
rect 1548 92491 1554 92543
rect 894 92371 1554 92491
rect 894 92319 900 92371
rect 1548 92319 1554 92371
rect 894 92199 1554 92319
rect 894 92147 900 92199
rect 1548 92147 1554 92199
rect 894 92027 1554 92147
rect 894 91975 900 92027
rect 1548 91975 1554 92027
rect 894 91855 1554 91975
rect 894 91803 900 91855
rect 1548 91803 1554 91855
rect 894 91683 1554 91803
rect 894 91631 900 91683
rect 1548 91631 1554 91683
rect 894 91511 1554 91631
rect 894 91459 900 91511
rect 1548 91459 1554 91511
rect 894 91339 1554 91459
rect 894 91287 900 91339
rect 1548 91287 1554 91339
rect 894 91167 1554 91287
rect 894 91115 900 91167
rect 1548 91115 1554 91167
rect 894 90995 1554 91115
rect 894 90943 900 90995
rect 1548 90943 1554 90995
rect 894 90823 1554 90943
rect 894 90771 900 90823
rect 1548 90771 1554 90823
rect 894 90651 1554 90771
rect 894 90599 900 90651
rect 1548 90599 1554 90651
rect 894 90479 1554 90599
rect 894 90427 900 90479
rect 1548 90427 1554 90479
rect 894 90307 1554 90427
rect 894 90255 900 90307
rect 1548 90255 1554 90307
rect 894 90135 1554 90255
rect 894 90083 900 90135
rect 1548 90083 1554 90135
rect 894 89963 1554 90083
rect 894 89911 900 89963
rect 1548 89911 1554 89963
rect 894 89791 1554 89911
rect 894 89739 900 89791
rect 1548 89739 1554 89791
rect 894 89619 1554 89739
rect 894 89567 900 89619
rect 1548 89567 1554 89619
rect 894 89447 1554 89567
rect 894 89395 900 89447
rect 1548 89395 1554 89447
rect 894 89275 1554 89395
rect 894 89223 900 89275
rect 1548 89223 1554 89275
rect 894 89103 1554 89223
rect 894 89051 900 89103
rect 1548 89051 1554 89103
rect 894 88931 1554 89051
rect 894 88879 900 88931
rect 1548 88879 1554 88931
rect 894 88759 1554 88879
rect 894 88707 900 88759
rect 1548 88707 1554 88759
rect 894 88587 1554 88707
rect 894 88535 900 88587
rect 1548 88535 1554 88587
rect 894 88415 1554 88535
rect 894 88363 900 88415
rect 1548 88363 1554 88415
rect 894 88243 1554 88363
rect 894 88191 900 88243
rect 1548 88191 1554 88243
rect 894 88071 1554 88191
rect 894 88019 900 88071
rect 1548 88019 1554 88071
rect 894 87899 1554 88019
rect 894 87847 900 87899
rect 1548 87847 1554 87899
rect 894 87727 1554 87847
rect 894 87675 900 87727
rect 1548 87675 1554 87727
rect 894 87555 1554 87675
rect 894 87503 900 87555
rect 1548 87503 1554 87555
rect 894 87383 1554 87503
rect 894 87331 900 87383
rect 1548 87331 1554 87383
rect 894 87211 1554 87331
rect 894 87159 900 87211
rect 1548 87159 1554 87211
rect 894 87039 1554 87159
rect 894 86987 900 87039
rect 1548 86987 1554 87039
rect 894 86867 1554 86987
rect 894 86815 900 86867
rect 1548 86815 1554 86867
rect 894 86695 1554 86815
rect 894 86643 900 86695
rect 1548 86643 1554 86695
rect 894 86523 1554 86643
rect 894 86471 900 86523
rect 1548 86471 1554 86523
rect 894 86351 1554 86471
rect 894 86299 900 86351
rect 1548 86299 1554 86351
rect 894 86179 1554 86299
rect 894 86127 900 86179
rect 1548 86127 1554 86179
rect 894 86007 1554 86127
rect 894 85955 900 86007
rect 1548 85955 1554 86007
rect 894 85835 1554 85955
rect 894 85783 900 85835
rect 1548 85783 1554 85835
rect 894 85663 1554 85783
rect 894 85611 900 85663
rect 1548 85611 1554 85663
rect 894 85491 1554 85611
rect 894 85439 900 85491
rect 1548 85439 1554 85491
rect 894 85319 1554 85439
rect 894 85267 900 85319
rect 1548 85267 1554 85319
rect 894 85147 1554 85267
rect 894 85095 900 85147
rect 1548 85095 1554 85147
rect 894 84975 1554 85095
rect 894 84923 900 84975
rect 1548 84923 1554 84975
rect 894 84803 1554 84923
rect 894 84751 900 84803
rect 1548 84751 1554 84803
rect 894 84631 1554 84751
rect 894 84579 900 84631
rect 1548 84579 1554 84631
rect 894 84459 1554 84579
rect 894 84407 900 84459
rect 1548 84407 1554 84459
rect 894 84287 1554 84407
rect 894 84235 900 84287
rect 1548 84235 1554 84287
rect 894 84115 1554 84235
rect 894 84063 900 84115
rect 1548 84063 1554 84115
rect 894 83943 1554 84063
rect 894 83891 900 83943
rect 1548 83891 1554 83943
rect 894 83771 1554 83891
rect 894 83719 900 83771
rect 1548 83719 1554 83771
rect 894 83599 1554 83719
rect 894 83547 900 83599
rect 1548 83547 1554 83599
rect 894 83427 1554 83547
rect 894 83375 900 83427
rect 1548 83375 1554 83427
rect 894 83255 1554 83375
rect 894 83203 900 83255
rect 1548 83203 1554 83255
rect 894 83083 1554 83203
rect 894 83031 900 83083
rect 1548 83031 1554 83083
rect 894 82911 1554 83031
rect 894 82859 900 82911
rect 1548 82859 1554 82911
rect 894 82739 1554 82859
rect 894 82687 900 82739
rect 1548 82687 1554 82739
rect 894 82567 1554 82687
rect 894 82515 900 82567
rect 1548 82515 1554 82567
rect 894 82395 1554 82515
rect 894 82343 900 82395
rect 1548 82343 1554 82395
rect 894 82223 1554 82343
rect 894 82171 900 82223
rect 1548 82171 1554 82223
rect 894 82051 1554 82171
rect 894 81999 900 82051
rect 1548 81999 1554 82051
rect 894 81879 1554 81999
rect 894 81827 900 81879
rect 1548 81827 1554 81879
rect 894 81707 1554 81827
rect 894 81655 900 81707
rect 1548 81655 1554 81707
rect 894 81535 1554 81655
rect 894 81483 900 81535
rect 1548 81483 1554 81535
rect 894 81363 1554 81483
rect 894 81311 900 81363
rect 1548 81311 1554 81363
rect 894 81191 1554 81311
rect 894 81139 900 81191
rect 1548 81139 1554 81191
rect 894 81019 1554 81139
rect 894 80967 900 81019
rect 1548 80967 1554 81019
rect 894 80847 1554 80967
rect 894 80795 900 80847
rect 1548 80795 1554 80847
rect 894 80675 1554 80795
rect 894 80623 900 80675
rect 1548 80623 1554 80675
rect 894 80503 1554 80623
rect 894 80451 900 80503
rect 1548 80451 1554 80503
rect 894 80331 1554 80451
rect 894 80279 900 80331
rect 1548 80279 1554 80331
rect 894 80159 1554 80279
rect 894 80107 900 80159
rect 1548 80107 1554 80159
rect 894 79987 1554 80107
rect 894 79935 900 79987
rect 1548 79935 1554 79987
rect 894 79815 1554 79935
rect 894 79763 900 79815
rect 1548 79763 1554 79815
rect 894 79643 1554 79763
rect 894 79591 900 79643
rect 1548 79591 1554 79643
rect 894 79471 1554 79591
rect 894 79419 900 79471
rect 1548 79419 1554 79471
rect 894 79299 1554 79419
rect 894 79247 900 79299
rect 1548 79247 1554 79299
rect 894 79127 1554 79247
rect 894 79075 900 79127
rect 1548 79075 1554 79127
rect 894 78955 1554 79075
rect 894 78903 900 78955
rect 1548 78903 1554 78955
rect 894 78783 1554 78903
rect 894 78731 900 78783
rect 1548 78731 1554 78783
rect 894 78611 1554 78731
rect 894 78559 900 78611
rect 1548 78559 1554 78611
rect 894 78439 1554 78559
rect 894 78387 900 78439
rect 1548 78387 1554 78439
rect 894 78267 1554 78387
rect 894 78215 900 78267
rect 1548 78215 1554 78267
rect 894 78095 1554 78215
rect 894 78043 900 78095
rect 1548 78043 1554 78095
rect 894 77923 1554 78043
rect 894 77871 900 77923
rect 1548 77871 1554 77923
rect 894 77751 1554 77871
rect 894 77699 900 77751
rect 1548 77699 1554 77751
rect 894 77579 1554 77699
rect 894 77527 900 77579
rect 1548 77527 1554 77579
rect 894 77407 1554 77527
rect 894 77355 900 77407
rect 1548 77355 1554 77407
rect 894 77235 1554 77355
rect 894 77183 900 77235
rect 1548 77183 1554 77235
rect 894 77063 1554 77183
rect 894 77011 900 77063
rect 1548 77011 1554 77063
rect 894 76891 1554 77011
rect 894 76839 900 76891
rect 1548 76839 1554 76891
rect 894 76719 1554 76839
rect 894 76667 900 76719
rect 1548 76667 1554 76719
rect 894 76547 1554 76667
rect 894 76495 900 76547
rect 1548 76495 1554 76547
rect 894 76375 1554 76495
rect 894 76323 900 76375
rect 1548 76323 1554 76375
rect 894 76203 1554 76323
rect 894 76151 900 76203
rect 1548 76151 1554 76203
rect 894 76031 1554 76151
rect 894 75979 900 76031
rect 1548 75979 1554 76031
rect 894 75859 1554 75979
rect 894 75807 900 75859
rect 1548 75807 1554 75859
rect 894 75687 1554 75807
rect 894 75635 900 75687
rect 1548 75635 1554 75687
rect 894 75515 1554 75635
rect 894 75463 900 75515
rect 1548 75463 1554 75515
rect 894 75343 1554 75463
rect 894 75291 900 75343
rect 1548 75291 1554 75343
rect 894 75171 1554 75291
rect 894 75119 900 75171
rect 1548 75119 1554 75171
rect 894 74999 1554 75119
rect 894 74947 900 74999
rect 1548 74947 1554 74999
rect 894 74827 1554 74947
rect 894 74775 900 74827
rect 1548 74775 1554 74827
rect 894 74655 1554 74775
rect 894 74603 900 74655
rect 1548 74603 1554 74655
rect 894 74483 1554 74603
rect 894 74431 900 74483
rect 1548 74431 1554 74483
rect 894 74311 1554 74431
rect 894 74259 900 74311
rect 1548 74259 1554 74311
rect 894 74139 1554 74259
rect 894 74087 900 74139
rect 1548 74087 1554 74139
rect 894 73967 1554 74087
rect 894 73915 900 73967
rect 1548 73915 1554 73967
rect 894 73795 1554 73915
rect 894 73743 900 73795
rect 1548 73743 1554 73795
rect 894 73623 1554 73743
rect 894 73571 900 73623
rect 1548 73571 1554 73623
rect 894 73451 1554 73571
rect 894 73399 900 73451
rect 1548 73399 1554 73451
rect 894 73279 1554 73399
rect 894 73227 900 73279
rect 1548 73227 1554 73279
rect 894 73107 1554 73227
rect 894 73055 900 73107
rect 1548 73055 1554 73107
rect 894 72935 1554 73055
rect 894 72883 900 72935
rect 1548 72883 1554 72935
rect 894 72763 1554 72883
rect 894 72711 900 72763
rect 1548 72711 1554 72763
rect 894 72591 1554 72711
rect 894 72539 900 72591
rect 1548 72539 1554 72591
rect 894 72419 1554 72539
rect 894 72367 900 72419
rect 1548 72367 1554 72419
rect 894 72247 1554 72367
rect 894 72195 900 72247
rect 1548 72195 1554 72247
rect 894 72075 1554 72195
rect 894 72023 900 72075
rect 1548 72023 1554 72075
rect 894 71903 1554 72023
rect 894 71851 900 71903
rect 1548 71851 1554 71903
rect 894 71731 1554 71851
rect 894 71679 900 71731
rect 1548 71679 1554 71731
rect 894 71559 1554 71679
rect 894 71507 900 71559
rect 1548 71507 1554 71559
rect 894 71387 1554 71507
rect 894 71335 900 71387
rect 1548 71335 1554 71387
rect 894 71215 1554 71335
rect 894 71163 900 71215
rect 1548 71163 1554 71215
rect 894 71043 1554 71163
rect 894 70991 900 71043
rect 1548 70991 1554 71043
rect 894 70871 1554 70991
rect 894 70819 900 70871
rect 1548 70819 1554 70871
rect 894 70699 1554 70819
rect 894 70647 900 70699
rect 1548 70647 1554 70699
rect 894 70527 1554 70647
rect 894 70475 900 70527
rect 1548 70475 1554 70527
rect 894 70355 1554 70475
rect 894 70303 900 70355
rect 1548 70303 1554 70355
rect 894 70183 1554 70303
rect 894 70131 900 70183
rect 1548 70131 1554 70183
rect 894 70011 1554 70131
rect 894 69959 900 70011
rect 1548 69959 1554 70011
rect 894 69839 1554 69959
rect 894 69787 900 69839
rect 1548 69787 1554 69839
rect 894 69667 1554 69787
rect 894 69615 900 69667
rect 1548 69615 1554 69667
rect 894 69495 1554 69615
rect 894 69443 900 69495
rect 1548 69443 1554 69495
rect 894 69323 1554 69443
rect 894 69271 900 69323
rect 1548 69271 1554 69323
rect 894 69151 1554 69271
rect 894 69099 900 69151
rect 1548 69099 1554 69151
rect 894 68979 1554 69099
rect 894 68927 900 68979
rect 1548 68927 1554 68979
rect 894 68807 1554 68927
rect 894 68755 900 68807
rect 1548 68755 1554 68807
rect 894 68635 1554 68755
rect 894 68583 900 68635
rect 1548 68583 1554 68635
rect 894 68463 1554 68583
rect 894 68411 900 68463
rect 1548 68411 1554 68463
rect 894 68291 1554 68411
rect 894 68239 900 68291
rect 1548 68239 1554 68291
rect 894 68119 1554 68239
rect 894 68067 900 68119
rect 1548 68067 1554 68119
rect 894 67947 1554 68067
rect 894 67895 900 67947
rect 1548 67895 1554 67947
rect 894 67775 1554 67895
rect 894 67723 900 67775
rect 1548 67723 1554 67775
rect 894 67603 1554 67723
rect 894 67551 900 67603
rect 1548 67551 1554 67603
rect 894 67431 1554 67551
rect 894 67379 900 67431
rect 1548 67379 1554 67431
rect 894 67259 1554 67379
rect 894 67207 900 67259
rect 1548 67207 1554 67259
rect 894 67087 1554 67207
rect 894 67035 900 67087
rect 1548 67035 1554 67087
rect 894 66915 1554 67035
rect 894 66863 900 66915
rect 1548 66863 1554 66915
rect 894 66743 1554 66863
rect 894 66691 900 66743
rect 1548 66691 1554 66743
rect 894 66571 1554 66691
rect 894 66519 900 66571
rect 1548 66519 1554 66571
rect 894 66399 1554 66519
rect 894 66347 900 66399
rect 1548 66347 1554 66399
rect 894 66227 1554 66347
rect 894 66175 900 66227
rect 1548 66175 1554 66227
rect 894 66055 1554 66175
rect 894 66003 900 66055
rect 1548 66003 1554 66055
rect 894 65883 1554 66003
rect 894 65831 900 65883
rect 1548 65831 1554 65883
rect 894 65711 1554 65831
rect 894 65659 900 65711
rect 1548 65659 1554 65711
rect 894 65539 1554 65659
rect 894 65487 900 65539
rect 1548 65487 1554 65539
rect 894 65367 1554 65487
rect 894 65315 900 65367
rect 1548 65315 1554 65367
rect 894 65195 1554 65315
rect 894 65143 900 65195
rect 1548 65143 1554 65195
rect 894 65023 1554 65143
rect 894 64971 900 65023
rect 1548 64971 1554 65023
rect 894 64851 1554 64971
rect 894 64799 900 64851
rect 1548 64799 1554 64851
rect 894 64679 1554 64799
rect 894 64627 900 64679
rect 1548 64627 1554 64679
rect 894 64507 1554 64627
rect 894 64455 900 64507
rect 1548 64455 1554 64507
rect 894 64335 1554 64455
rect 894 64283 900 64335
rect 1548 64283 1554 64335
rect 894 64163 1554 64283
rect 894 64111 900 64163
rect 1548 64111 1554 64163
rect 894 63991 1554 64111
rect 894 63939 900 63991
rect 1548 63939 1554 63991
rect 894 63819 1554 63939
rect 894 63767 900 63819
rect 1548 63767 1554 63819
rect 894 63647 1554 63767
rect 894 63595 900 63647
rect 1548 63595 1554 63647
rect 894 63475 1554 63595
rect 894 63423 900 63475
rect 1548 63423 1554 63475
rect 894 63303 1554 63423
rect 894 63251 900 63303
rect 1548 63251 1554 63303
rect 894 63131 1554 63251
rect 894 63079 900 63131
rect 1548 63079 1554 63131
rect 894 62959 1554 63079
rect 894 62907 900 62959
rect 1548 62907 1554 62959
rect 894 62787 1554 62907
rect 894 62735 900 62787
rect 1548 62735 1554 62787
rect 894 62615 1554 62735
rect 894 62563 900 62615
rect 1548 62563 1554 62615
rect 894 62443 1554 62563
rect 894 62391 900 62443
rect 1548 62391 1554 62443
rect 894 62271 1554 62391
rect 894 62219 900 62271
rect 1548 62219 1554 62271
rect 894 62099 1554 62219
rect 894 62047 900 62099
rect 1548 62047 1554 62099
rect 894 61927 1554 62047
rect 894 61875 900 61927
rect 1548 61875 1554 61927
rect 894 61755 1554 61875
rect 894 61703 900 61755
rect 1548 61703 1554 61755
rect 894 61583 1554 61703
rect 894 61531 900 61583
rect 1548 61531 1554 61583
rect 894 61411 1554 61531
rect 894 61359 900 61411
rect 1548 61359 1554 61411
rect 894 61239 1554 61359
rect 894 61187 900 61239
rect 1548 61187 1554 61239
rect 894 61067 1554 61187
rect 894 61015 900 61067
rect 1548 61015 1554 61067
rect 894 60895 1554 61015
rect 894 60843 900 60895
rect 1548 60843 1554 60895
rect 894 60723 1554 60843
rect 894 60671 900 60723
rect 1548 60671 1554 60723
rect 894 60551 1554 60671
rect 894 60499 900 60551
rect 1548 60499 1554 60551
rect 894 60379 1554 60499
rect 894 60327 900 60379
rect 1548 60327 1554 60379
rect 894 60207 1554 60327
rect 894 60155 900 60207
rect 1548 60155 1554 60207
rect 894 60035 1554 60155
rect 894 59983 900 60035
rect 1548 59983 1554 60035
rect 894 59863 1554 59983
rect 894 59811 900 59863
rect 1548 59811 1554 59863
rect 894 59691 1554 59811
rect 894 59639 900 59691
rect 1548 59639 1554 59691
rect 894 59519 1554 59639
rect 894 59467 900 59519
rect 1548 59467 1554 59519
rect 894 59347 1554 59467
rect 894 59295 900 59347
rect 1548 59295 1554 59347
rect 894 59175 1554 59295
rect 894 59123 900 59175
rect 1548 59123 1554 59175
rect 894 59003 1554 59123
rect 894 58951 900 59003
rect 1548 58951 1554 59003
rect 894 58831 1554 58951
rect 894 58779 900 58831
rect 1548 58779 1554 58831
rect 894 58659 1554 58779
rect 894 58607 900 58659
rect 1548 58607 1554 58659
rect 894 58487 1554 58607
rect 894 58435 900 58487
rect 1548 58435 1554 58487
rect 894 58315 1554 58435
rect 894 58263 900 58315
rect 1548 58263 1554 58315
rect 894 58143 1554 58263
rect 894 58091 900 58143
rect 1548 58091 1554 58143
rect 894 57971 1554 58091
rect 894 57919 900 57971
rect 1548 57919 1554 57971
rect 894 57799 1554 57919
rect 894 57747 900 57799
rect 1548 57747 1554 57799
rect 894 57627 1554 57747
rect 894 57575 900 57627
rect 1548 57575 1554 57627
rect 894 57455 1554 57575
rect 894 57403 900 57455
rect 1548 57403 1554 57455
rect 894 57283 1554 57403
rect 894 57231 900 57283
rect 1548 57231 1554 57283
rect 894 57111 1554 57231
rect 894 57059 900 57111
rect 1548 57059 1554 57111
rect 894 56939 1554 57059
rect 894 56887 900 56939
rect 1548 56887 1554 56939
rect 894 56767 1554 56887
rect 894 56715 900 56767
rect 1548 56715 1554 56767
rect 894 56595 1554 56715
rect 894 56543 900 56595
rect 1548 56543 1554 56595
rect 894 56423 1554 56543
rect 894 56371 900 56423
rect 1548 56371 1554 56423
rect 894 56251 1554 56371
rect 894 56199 900 56251
rect 1548 56199 1554 56251
rect 894 56079 1554 56199
rect 894 56027 900 56079
rect 1548 56027 1554 56079
rect 894 55907 1554 56027
rect 894 55855 900 55907
rect 1548 55855 1554 55907
rect 894 55735 1554 55855
rect 894 55683 900 55735
rect 1548 55683 1554 55735
rect 894 55563 1554 55683
rect 894 55511 900 55563
rect 1548 55511 1554 55563
rect 894 55391 1554 55511
rect 894 55339 900 55391
rect 1548 55339 1554 55391
rect 894 55219 1554 55339
rect 894 55167 900 55219
rect 1548 55167 1554 55219
rect 894 55047 1554 55167
rect 894 54995 900 55047
rect 1548 54995 1554 55047
rect 894 54875 1554 54995
rect 894 54823 900 54875
rect 1548 54823 1554 54875
rect 894 54703 1554 54823
rect 894 54651 900 54703
rect 1548 54651 1554 54703
rect 894 54531 1554 54651
rect 894 54479 900 54531
rect 1548 54479 1554 54531
rect 894 54359 1554 54479
rect 894 54307 900 54359
rect 1548 54307 1554 54359
rect 894 54187 1554 54307
rect 894 54135 900 54187
rect 1548 54135 1554 54187
rect 894 54015 1554 54135
rect 894 53963 900 54015
rect 1548 53963 1554 54015
rect 894 53843 1554 53963
rect 894 53791 900 53843
rect 1548 53791 1554 53843
rect 894 53671 1554 53791
rect 894 53619 900 53671
rect 1548 53619 1554 53671
rect 894 53499 1554 53619
rect 894 53447 900 53499
rect 1548 53447 1554 53499
rect 894 53327 1554 53447
rect 894 53275 900 53327
rect 1548 53275 1554 53327
rect 894 53155 1554 53275
rect 894 53103 900 53155
rect 1548 53103 1554 53155
rect 894 52983 1554 53103
rect 894 52931 900 52983
rect 1548 52931 1554 52983
rect 894 52811 1554 52931
rect 894 52759 900 52811
rect 1548 52759 1554 52811
rect 894 52639 1554 52759
rect 894 52587 900 52639
rect 1548 52587 1554 52639
rect 894 52467 1554 52587
rect 894 52415 900 52467
rect 1548 52415 1554 52467
rect 894 52295 1554 52415
rect 894 52243 900 52295
rect 1548 52243 1554 52295
rect 894 52123 1554 52243
rect 894 52071 900 52123
rect 1548 52071 1554 52123
rect 894 51951 1554 52071
rect 894 51899 900 51951
rect 1548 51899 1554 51951
rect 894 51779 1554 51899
rect 894 51727 900 51779
rect 1548 51727 1554 51779
rect 894 51607 1554 51727
rect 894 51555 900 51607
rect 1548 51555 1554 51607
rect 894 51435 1554 51555
rect 894 51383 900 51435
rect 1548 51383 1554 51435
rect 894 51263 1554 51383
rect 894 51211 900 51263
rect 1548 51211 1554 51263
rect 894 51091 1554 51211
rect 894 51039 900 51091
rect 1548 51039 1554 51091
rect 894 50919 1554 51039
rect 894 50867 900 50919
rect 1548 50867 1554 50919
rect 894 50747 1554 50867
rect 894 50695 900 50747
rect 1548 50695 1554 50747
rect 894 50575 1554 50695
rect 894 50523 900 50575
rect 1548 50523 1554 50575
rect 894 50403 1554 50523
rect 894 50351 900 50403
rect 1548 50351 1554 50403
rect 894 50231 1554 50351
rect 894 50179 900 50231
rect 1548 50179 1554 50231
rect 894 50059 1554 50179
rect 894 50007 900 50059
rect 1548 50007 1554 50059
rect 894 49887 1554 50007
rect 894 49835 900 49887
rect 1548 49835 1554 49887
rect 894 49715 1554 49835
rect 894 49663 900 49715
rect 1548 49663 1554 49715
rect 894 49543 1554 49663
rect 894 49491 900 49543
rect 1548 49491 1554 49543
rect 894 49371 1554 49491
rect 894 49319 900 49371
rect 1548 49319 1554 49371
rect 894 49199 1554 49319
rect 894 49147 900 49199
rect 1548 49147 1554 49199
rect 894 49027 1554 49147
rect 894 48975 900 49027
rect 1548 48975 1554 49027
rect 894 48855 1554 48975
rect 894 48803 900 48855
rect 1548 48803 1554 48855
rect 894 48683 1554 48803
rect 894 48631 900 48683
rect 1548 48631 1554 48683
rect 894 48511 1554 48631
rect 894 48459 900 48511
rect 1548 48459 1554 48511
rect 894 48339 1554 48459
rect 894 48287 900 48339
rect 1548 48287 1554 48339
rect 894 48167 1554 48287
rect 894 48115 900 48167
rect 1548 48115 1554 48167
rect 894 47995 1554 48115
rect 894 47943 900 47995
rect 1548 47943 1554 47995
rect 894 47823 1554 47943
rect 894 47771 900 47823
rect 1548 47771 1554 47823
rect 894 47651 1554 47771
rect 894 47599 900 47651
rect 1548 47599 1554 47651
rect 894 47479 1554 47599
rect 894 47427 900 47479
rect 1548 47427 1554 47479
rect 894 47307 1554 47427
rect 894 47255 900 47307
rect 1548 47255 1554 47307
rect 894 47135 1554 47255
rect 894 47083 900 47135
rect 1548 47083 1554 47135
rect 894 46963 1554 47083
rect 894 46911 900 46963
rect 1548 46911 1554 46963
rect 894 46791 1554 46911
rect 894 46739 900 46791
rect 1548 46739 1554 46791
rect 894 46619 1554 46739
rect 894 46567 900 46619
rect 1548 46567 1554 46619
rect 894 46447 1554 46567
rect 894 46395 900 46447
rect 1548 46395 1554 46447
rect 894 46275 1554 46395
rect 894 46223 900 46275
rect 1548 46223 1554 46275
rect 894 46103 1554 46223
rect 894 46051 900 46103
rect 1548 46051 1554 46103
rect 894 45931 1554 46051
rect 894 45879 900 45931
rect 1548 45879 1554 45931
rect 894 45759 1554 45879
rect 894 45707 900 45759
rect 1548 45707 1554 45759
rect 894 45587 1554 45707
rect 894 45535 900 45587
rect 1548 45535 1554 45587
rect 894 45415 1554 45535
rect 894 45363 900 45415
rect 1548 45363 1554 45415
rect 894 45243 1554 45363
rect 894 45191 900 45243
rect 1548 45191 1554 45243
rect 894 45071 1554 45191
rect 894 45019 900 45071
rect 1548 45019 1554 45071
rect 894 44899 1554 45019
rect 894 44847 900 44899
rect 1548 44847 1554 44899
rect 894 44727 1554 44847
rect 894 44675 900 44727
rect 1548 44675 1554 44727
rect 894 44555 1554 44675
rect 894 44503 900 44555
rect 1548 44503 1554 44555
rect 894 44383 1554 44503
rect 894 44331 900 44383
rect 1548 44331 1554 44383
rect 894 44211 1554 44331
rect 894 44159 900 44211
rect 1548 44159 1554 44211
rect 894 44039 1554 44159
rect 894 43987 900 44039
rect 1548 43987 1554 44039
rect 894 43867 1554 43987
rect 894 43815 900 43867
rect 1548 43815 1554 43867
rect 894 43695 1554 43815
rect 894 43643 900 43695
rect 1548 43643 1554 43695
rect 894 43523 1554 43643
rect 894 43471 900 43523
rect 1548 43471 1554 43523
rect 894 43351 1554 43471
rect 894 43299 900 43351
rect 1548 43299 1554 43351
rect 894 43179 1554 43299
rect 894 43127 900 43179
rect 1548 43127 1554 43179
rect 894 43007 1554 43127
rect 894 42955 900 43007
rect 1548 42955 1554 43007
rect 894 42835 1554 42955
rect 894 42783 900 42835
rect 1548 42783 1554 42835
rect 894 42663 1554 42783
rect 894 42611 900 42663
rect 1548 42611 1554 42663
rect 894 42491 1554 42611
rect 894 42439 900 42491
rect 1548 42439 1554 42491
rect 894 42319 1554 42439
rect 894 42267 900 42319
rect 1548 42267 1554 42319
rect 894 42147 1554 42267
rect 894 42095 900 42147
rect 1548 42095 1554 42147
rect 894 41975 1554 42095
rect 894 41923 900 41975
rect 1548 41923 1554 41975
rect 894 41803 1554 41923
rect 894 41751 900 41803
rect 1548 41751 1554 41803
rect 894 41631 1554 41751
rect 894 41579 900 41631
rect 1548 41579 1554 41631
rect 894 41459 1554 41579
rect 894 41407 900 41459
rect 1548 41407 1554 41459
rect 894 41287 1554 41407
rect 894 41235 900 41287
rect 1548 41235 1554 41287
rect 894 41115 1554 41235
rect 894 41063 900 41115
rect 1548 41063 1554 41115
rect 894 40943 1554 41063
rect 894 40891 900 40943
rect 1548 40891 1554 40943
rect 894 40771 1554 40891
rect 894 40719 900 40771
rect 1548 40719 1554 40771
rect 894 40599 1554 40719
rect 894 40547 900 40599
rect 1548 40547 1554 40599
rect 894 40427 1554 40547
rect 894 40375 900 40427
rect 1548 40375 1554 40427
rect 894 40255 1554 40375
rect 894 40203 900 40255
rect 1548 40203 1554 40255
rect 894 40083 1554 40203
rect 894 40031 900 40083
rect 1548 40031 1554 40083
rect 894 39911 1554 40031
rect 894 39859 900 39911
rect 1548 39859 1554 39911
rect 894 39739 1554 39859
rect 894 39687 900 39739
rect 1548 39687 1554 39739
rect 894 39567 1554 39687
rect 894 39515 900 39567
rect 1548 39515 1554 39567
rect 894 39395 1554 39515
rect 894 39343 900 39395
rect 1548 39343 1554 39395
rect 894 39223 1554 39343
rect 894 39171 900 39223
rect 1548 39171 1554 39223
rect 894 39051 1554 39171
rect 894 38999 900 39051
rect 1548 38999 1554 39051
rect 894 38879 1554 38999
rect 894 38827 900 38879
rect 1548 38827 1554 38879
rect 894 38707 1554 38827
rect 894 38655 900 38707
rect 1548 38655 1554 38707
rect 894 38535 1554 38655
rect 894 38483 900 38535
rect 1548 38483 1554 38535
rect 894 38363 1554 38483
rect 894 38311 900 38363
rect 1548 38311 1554 38363
rect 894 38191 1554 38311
rect 894 38139 900 38191
rect 1548 38139 1554 38191
rect 894 38019 1554 38139
rect 894 37967 900 38019
rect 1548 37967 1554 38019
rect 894 37847 1554 37967
rect 894 37795 900 37847
rect 1548 37795 1554 37847
rect 894 37675 1554 37795
rect 894 37623 900 37675
rect 1548 37623 1554 37675
rect 894 37503 1554 37623
rect 894 37451 900 37503
rect 1548 37451 1554 37503
rect 894 37331 1554 37451
rect 894 37279 900 37331
rect 1548 37279 1554 37331
rect 894 37159 1554 37279
rect 894 37107 900 37159
rect 1548 37107 1554 37159
rect 894 36987 1554 37107
rect 894 36935 900 36987
rect 1548 36935 1554 36987
rect 894 36815 1554 36935
rect 894 36763 900 36815
rect 1548 36763 1554 36815
rect 894 36643 1554 36763
rect 894 36591 900 36643
rect 1548 36591 1554 36643
rect 894 36471 1554 36591
rect 894 36419 900 36471
rect 1548 36419 1554 36471
rect 894 36299 1554 36419
rect 894 36247 900 36299
rect 1548 36247 1554 36299
rect 894 36127 1554 36247
rect 894 36075 900 36127
rect 1548 36075 1554 36127
rect 894 35955 1554 36075
rect 894 35903 900 35955
rect 1548 35903 1554 35955
rect 894 35783 1554 35903
rect 894 35731 900 35783
rect 1548 35731 1554 35783
rect 894 35611 1554 35731
rect 894 35559 900 35611
rect 1548 35559 1554 35611
rect 894 35439 1554 35559
rect 894 35387 900 35439
rect 1548 35387 1554 35439
rect 894 35267 1554 35387
rect 894 35215 900 35267
rect 1548 35215 1554 35267
rect 894 35095 1554 35215
rect 894 35043 900 35095
rect 1548 35043 1554 35095
rect 894 34923 1554 35043
rect 894 34871 900 34923
rect 1548 34871 1554 34923
rect 894 34751 1554 34871
rect 894 34699 900 34751
rect 1548 34699 1554 34751
rect 894 34579 1554 34699
rect 894 34527 900 34579
rect 1548 34527 1554 34579
rect 894 34407 1554 34527
rect 894 34355 900 34407
rect 1548 34355 1554 34407
rect 894 34235 1554 34355
rect 894 34183 900 34235
rect 1548 34183 1554 34235
rect 894 34063 1554 34183
rect 894 34011 900 34063
rect 1548 34011 1554 34063
rect 894 33891 1554 34011
rect 894 33839 900 33891
rect 1548 33839 1554 33891
rect 894 33719 1554 33839
rect 894 33667 900 33719
rect 1548 33667 1554 33719
rect 894 33547 1554 33667
rect 894 33495 900 33547
rect 1548 33495 1554 33547
rect 894 33375 1554 33495
rect 894 33323 900 33375
rect 1548 33323 1554 33375
rect 894 33203 1554 33323
rect 894 33151 900 33203
rect 1548 33151 1554 33203
rect 894 33031 1554 33151
rect 894 32979 900 33031
rect 1548 32979 1554 33031
rect 894 32859 1554 32979
rect 894 32807 900 32859
rect 1548 32807 1554 32859
rect 894 32687 1554 32807
rect 894 32635 900 32687
rect 1548 32635 1554 32687
rect 894 32515 1554 32635
rect 894 32463 900 32515
rect 1548 32463 1554 32515
rect 894 32343 1554 32463
rect 894 32291 900 32343
rect 1548 32291 1554 32343
rect 894 32171 1554 32291
rect 894 32119 900 32171
rect 1548 32119 1554 32171
rect 894 31999 1554 32119
rect 894 31947 900 31999
rect 1548 31947 1554 31999
rect 894 31827 1554 31947
rect 894 31775 900 31827
rect 1548 31775 1554 31827
rect 894 31655 1554 31775
rect 894 31603 900 31655
rect 1548 31603 1554 31655
rect 894 31483 1554 31603
rect 894 31431 900 31483
rect 1548 31431 1554 31483
rect 894 31311 1554 31431
rect 894 31259 900 31311
rect 1548 31259 1554 31311
rect 894 31139 1554 31259
rect 894 31087 900 31139
rect 1548 31087 1554 31139
rect 894 30967 1554 31087
rect 894 30915 900 30967
rect 1548 30915 1554 30967
rect 894 30795 1554 30915
rect 894 30743 900 30795
rect 1548 30743 1554 30795
rect 894 30623 1554 30743
rect 894 30571 900 30623
rect 1548 30571 1554 30623
rect 894 30451 1554 30571
rect 894 30399 900 30451
rect 1548 30399 1554 30451
rect 894 30279 1554 30399
rect 894 30227 900 30279
rect 1548 30227 1554 30279
rect 894 30107 1554 30227
rect 894 30055 900 30107
rect 1548 30055 1554 30107
rect 894 29935 1554 30055
rect 894 29883 900 29935
rect 1548 29883 1554 29935
rect 894 29763 1554 29883
rect 894 29711 900 29763
rect 1548 29711 1554 29763
rect 894 29591 1554 29711
rect 894 29539 900 29591
rect 1548 29539 1554 29591
rect 894 29419 1554 29539
rect 894 29367 900 29419
rect 1548 29367 1554 29419
rect 894 29247 1554 29367
rect 894 29195 900 29247
rect 1548 29195 1554 29247
rect 894 29075 1554 29195
rect 894 29023 900 29075
rect 1548 29023 1554 29075
rect 894 28903 1554 29023
rect 894 28851 900 28903
rect 1548 28851 1554 28903
rect 894 28731 1554 28851
rect 894 28679 900 28731
rect 1548 28679 1554 28731
rect 894 28559 1554 28679
rect 894 28507 900 28559
rect 1548 28507 1554 28559
rect 894 28387 1554 28507
rect 894 28335 900 28387
rect 1548 28335 1554 28387
rect 894 28215 1554 28335
rect 894 28163 900 28215
rect 1548 28163 1554 28215
rect 894 28043 1554 28163
rect 894 27991 900 28043
rect 1548 27991 1554 28043
rect 894 27871 1554 27991
rect 894 27819 900 27871
rect 1548 27819 1554 27871
rect 894 27699 1554 27819
rect 894 27647 900 27699
rect 1548 27647 1554 27699
rect 894 27527 1554 27647
rect 894 27475 900 27527
rect 1548 27475 1554 27527
rect 894 27355 1554 27475
rect 894 27303 900 27355
rect 1548 27303 1554 27355
rect 894 27183 1554 27303
rect 894 27131 900 27183
rect 1548 27131 1554 27183
rect 894 27011 1554 27131
rect 894 26959 900 27011
rect 1548 26959 1554 27011
rect 894 26839 1554 26959
rect 894 26787 900 26839
rect 1548 26787 1554 26839
rect 894 26667 1554 26787
rect 894 26615 900 26667
rect 1548 26615 1554 26667
rect 894 26495 1554 26615
rect 894 26443 900 26495
rect 1548 26443 1554 26495
rect 894 26323 1554 26443
rect 894 26271 900 26323
rect 1548 26271 1554 26323
rect 894 26151 1554 26271
rect 894 26099 900 26151
rect 1548 26099 1554 26151
rect 894 25979 1554 26099
rect 894 25927 900 25979
rect 1548 25927 1554 25979
rect 894 25807 1554 25927
rect 894 25755 900 25807
rect 1548 25755 1554 25807
rect 894 25635 1554 25755
rect 894 25583 900 25635
rect 1548 25583 1554 25635
rect 894 25463 1554 25583
rect 894 25411 900 25463
rect 1548 25411 1554 25463
rect 894 25291 1554 25411
rect 894 25239 900 25291
rect 1548 25239 1554 25291
rect 894 25119 1554 25239
rect 894 25067 900 25119
rect 1548 25067 1554 25119
rect 894 24947 1554 25067
rect 894 24895 900 24947
rect 1548 24895 1554 24947
rect 894 24775 1554 24895
rect 894 24723 900 24775
rect 1548 24723 1554 24775
rect 894 24603 1554 24723
rect 894 24551 900 24603
rect 1548 24551 1554 24603
rect 894 24431 1554 24551
rect 894 24379 900 24431
rect 1548 24379 1554 24431
rect 894 24259 1554 24379
rect 894 24207 900 24259
rect 1548 24207 1554 24259
rect 894 24087 1554 24207
rect 894 24035 900 24087
rect 1548 24035 1554 24087
rect 894 23915 1554 24035
rect 894 23863 900 23915
rect 1548 23863 1554 23915
rect 894 23743 1554 23863
rect 894 23691 900 23743
rect 1548 23691 1554 23743
rect 894 23571 1554 23691
rect 894 23519 900 23571
rect 1548 23519 1554 23571
rect 894 23399 1554 23519
rect 894 23347 900 23399
rect 1548 23347 1554 23399
rect 894 23227 1554 23347
rect 894 23175 900 23227
rect 1548 23175 1554 23227
rect 894 23055 1554 23175
rect 894 23003 900 23055
rect 1548 23003 1554 23055
rect 894 22883 1554 23003
rect 894 22831 900 22883
rect 1548 22831 1554 22883
rect 894 22711 1554 22831
rect 894 22659 900 22711
rect 1548 22659 1554 22711
rect 894 22539 1554 22659
rect 894 22487 900 22539
rect 1548 22487 1554 22539
rect 894 22367 1554 22487
rect 894 22315 900 22367
rect 1548 22315 1554 22367
rect 894 22195 1554 22315
rect 894 22143 900 22195
rect 1548 22143 1554 22195
rect 894 22023 1554 22143
rect 894 21971 900 22023
rect 1548 21971 1554 22023
rect 894 21851 1554 21971
rect 894 21799 900 21851
rect 1548 21799 1554 21851
rect 894 21679 1554 21799
rect 894 21627 900 21679
rect 1548 21627 1554 21679
rect 894 21507 1554 21627
rect 894 21455 900 21507
rect 1548 21455 1554 21507
rect 894 21335 1554 21455
rect 894 21283 900 21335
rect 1548 21283 1554 21335
rect 894 21163 1554 21283
rect 894 21111 900 21163
rect 1548 21111 1554 21163
rect 894 20991 1554 21111
rect 894 20939 900 20991
rect 1548 20939 1554 20991
rect 894 20819 1554 20939
rect 894 20767 900 20819
rect 1548 20767 1554 20819
rect 894 20647 1554 20767
rect 894 20595 900 20647
rect 1548 20595 1554 20647
rect 894 20475 1554 20595
rect 894 20423 900 20475
rect 1548 20423 1554 20475
rect 894 20303 1554 20423
rect 894 20251 900 20303
rect 1548 20251 1554 20303
rect 894 20131 1554 20251
rect 894 20079 900 20131
rect 1548 20079 1554 20131
rect 894 19959 1554 20079
rect 894 19907 900 19959
rect 1548 19907 1554 19959
rect 894 19787 1554 19907
rect 894 19735 900 19787
rect 1548 19735 1554 19787
rect 894 19615 1554 19735
rect 894 19563 900 19615
rect 1548 19563 1554 19615
rect 894 19443 1554 19563
rect 894 19391 900 19443
rect 1548 19391 1554 19443
rect 894 19271 1554 19391
rect 894 19219 900 19271
rect 1548 19219 1554 19271
rect 894 19099 1554 19219
rect 894 19047 900 19099
rect 1548 19047 1554 19099
rect 894 18927 1554 19047
rect 894 18875 900 18927
rect 1548 18875 1554 18927
rect 894 18755 1554 18875
rect 894 18703 900 18755
rect 1548 18703 1554 18755
rect 894 18583 1554 18703
rect 894 18531 900 18583
rect 1548 18531 1554 18583
rect 894 18411 1554 18531
rect 894 18359 900 18411
rect 1548 18359 1554 18411
rect 894 18239 1554 18359
rect 894 18187 900 18239
rect 1548 18187 1554 18239
rect 894 18067 1554 18187
rect 894 18015 900 18067
rect 1548 18015 1554 18067
rect 894 17895 1554 18015
rect 894 17843 900 17895
rect 1548 17843 1554 17895
rect 894 17723 1554 17843
rect 894 17671 900 17723
rect 1548 17671 1554 17723
rect 894 17551 1554 17671
rect 894 17499 900 17551
rect 1548 17499 1554 17551
rect 894 17379 1554 17499
rect 894 17327 900 17379
rect 1548 17327 1554 17379
rect 894 17207 1554 17327
rect 894 17155 900 17207
rect 1548 17155 1554 17207
rect 894 17035 1554 17155
rect 894 16983 900 17035
rect 1548 16983 1554 17035
rect 894 16863 1554 16983
rect 894 16811 900 16863
rect 1548 16811 1554 16863
rect 894 16691 1554 16811
rect 894 16639 900 16691
rect 1548 16639 1554 16691
rect 894 16519 1554 16639
rect 894 16467 900 16519
rect 1548 16467 1554 16519
rect 894 16347 1554 16467
rect 894 16295 900 16347
rect 1548 16295 1554 16347
rect 894 16175 1554 16295
rect 894 16123 900 16175
rect 1548 16123 1554 16175
rect 894 16003 1554 16123
rect 894 15951 900 16003
rect 1548 15951 1554 16003
rect 894 15831 1554 15951
rect 894 15779 900 15831
rect 1548 15779 1554 15831
rect 894 15659 1554 15779
rect 894 15607 900 15659
rect 1548 15607 1554 15659
rect 894 15487 1554 15607
rect 894 15435 900 15487
rect 1548 15435 1554 15487
rect 894 15315 1554 15435
rect 894 15263 900 15315
rect 1548 15263 1554 15315
rect 894 15143 1554 15263
rect 894 15091 900 15143
rect 1548 15091 1554 15143
rect 894 14971 1554 15091
rect 894 14919 900 14971
rect 1548 14919 1554 14971
rect 894 14799 1554 14919
rect 894 14747 900 14799
rect 1548 14747 1554 14799
rect 894 14627 1554 14747
rect 894 14575 900 14627
rect 1548 14575 1554 14627
rect 894 14455 1554 14575
rect 894 14403 900 14455
rect 1548 14403 1554 14455
rect 894 14283 1554 14403
rect 894 14231 900 14283
rect 1548 14231 1554 14283
rect 894 14111 1554 14231
rect 894 14059 900 14111
rect 1548 14059 1554 14111
rect 894 13939 1554 14059
rect 894 13887 900 13939
rect 1548 13887 1554 13939
rect 894 13767 1554 13887
rect 894 13715 900 13767
rect 1548 13715 1554 13767
rect 894 13595 1554 13715
rect 894 13543 900 13595
rect 1548 13543 1554 13595
rect 894 13423 1554 13543
rect 894 13371 900 13423
rect 1548 13371 1554 13423
rect 894 13251 1554 13371
rect 894 13199 900 13251
rect 1548 13199 1554 13251
rect 894 13079 1554 13199
rect 894 13027 900 13079
rect 1548 13027 1554 13079
rect 894 12907 1554 13027
rect 894 12855 900 12907
rect 1548 12855 1554 12907
rect 894 12735 1554 12855
rect 894 12683 900 12735
rect 1548 12683 1554 12735
rect 894 12563 1554 12683
rect 894 12511 900 12563
rect 1548 12511 1554 12563
rect 894 12391 1554 12511
rect 894 12339 900 12391
rect 1548 12339 1554 12391
rect 894 12219 1554 12339
rect 894 12167 900 12219
rect 1548 12167 1554 12219
rect 894 12047 1554 12167
rect 894 11995 900 12047
rect 1548 11995 1554 12047
rect 894 11875 1554 11995
rect 894 11823 900 11875
rect 1548 11823 1554 11875
rect 894 11703 1554 11823
rect 894 11651 900 11703
rect 1548 11651 1554 11703
rect 894 11531 1554 11651
rect 894 11479 900 11531
rect 1548 11479 1554 11531
rect 894 11359 1554 11479
rect 894 11307 900 11359
rect 1548 11307 1554 11359
rect 894 11187 1554 11307
rect 894 11135 900 11187
rect 1548 11135 1554 11187
rect 894 11015 1554 11135
rect 894 10963 900 11015
rect 1548 10963 1554 11015
rect 894 10843 1554 10963
rect 894 10791 900 10843
rect 1548 10791 1554 10843
rect 894 10671 1554 10791
rect 894 10619 900 10671
rect 1548 10619 1554 10671
rect 894 10499 1554 10619
rect 894 10447 900 10499
rect 1548 10447 1554 10499
rect 894 10327 1554 10447
rect 894 10275 900 10327
rect 1548 10275 1554 10327
rect 894 10155 1554 10275
rect 894 10103 900 10155
rect 1548 10103 1554 10155
rect 894 9983 1554 10103
rect 894 9931 900 9983
rect 1548 9931 1554 9983
rect 894 9811 1554 9931
rect 894 9759 900 9811
rect 1548 9759 1554 9811
rect 894 9639 1554 9759
rect 894 9587 900 9639
rect 1548 9587 1554 9639
rect 894 9467 1554 9587
rect 894 9415 900 9467
rect 1548 9415 1554 9467
rect 894 9295 1554 9415
rect 894 9243 900 9295
rect 1548 9243 1554 9295
rect 894 9123 1554 9243
rect 894 9071 900 9123
rect 1548 9071 1554 9123
rect 894 8951 1554 9071
rect 894 8899 900 8951
rect 1548 8899 1554 8951
rect 894 8779 1554 8899
rect 894 8727 900 8779
rect 1548 8727 1554 8779
rect 894 8607 1554 8727
rect 894 8555 900 8607
rect 1548 8555 1554 8607
rect 894 8435 1554 8555
rect 894 8383 900 8435
rect 1548 8383 1554 8435
rect 894 8263 1554 8383
rect 894 8211 900 8263
rect 1548 8211 1554 8263
rect 894 8091 1554 8211
rect 894 8039 900 8091
rect 1548 8039 1554 8091
rect 894 7919 1554 8039
rect 894 7867 900 7919
rect 1548 7867 1554 7919
rect 894 7747 1554 7867
rect 894 7695 900 7747
rect 1548 7695 1554 7747
rect 894 7575 1554 7695
rect 894 7523 900 7575
rect 1548 7523 1554 7575
rect 894 7403 1554 7523
rect 894 7351 900 7403
rect 1548 7351 1554 7403
rect 894 7231 1554 7351
rect 894 7179 900 7231
rect 1548 7179 1554 7231
rect 894 7059 1554 7179
rect 894 7007 900 7059
rect 1548 7007 1554 7059
rect 894 6887 1554 7007
rect 894 6835 900 6887
rect 1548 6835 1554 6887
rect 894 6715 1554 6835
rect 894 6663 900 6715
rect 1548 6663 1554 6715
rect 894 6543 1554 6663
rect 894 6491 900 6543
rect 1548 6491 1554 6543
rect 894 6371 1554 6491
rect 894 6319 900 6371
rect 1548 6319 1554 6371
rect 894 6199 1554 6319
rect 894 6147 900 6199
rect 1548 6147 1554 6199
rect 894 6027 1554 6147
rect 894 5975 900 6027
rect 1548 5975 1554 6027
rect 894 5855 1554 5975
rect 894 5803 900 5855
rect 1548 5803 1554 5855
rect 894 5683 1554 5803
rect 894 5631 900 5683
rect 1548 5631 1554 5683
rect 894 5511 1554 5631
rect 894 5459 900 5511
rect 1548 5459 1554 5511
rect 894 5339 1554 5459
rect 894 5287 900 5339
rect 1548 5287 1554 5339
rect 894 5167 1554 5287
rect 894 5115 900 5167
rect 1548 5115 1554 5167
rect 894 4995 1554 5115
rect 894 4943 900 4995
rect 1548 4943 1554 4995
rect 894 4823 1554 4943
rect 894 4771 900 4823
rect 1548 4771 1554 4823
rect 894 4651 1554 4771
rect 894 4599 900 4651
rect 1548 4599 1554 4651
rect 894 4479 1554 4599
rect 894 4427 900 4479
rect 1548 4427 1554 4479
rect 894 4307 1554 4427
rect 894 4255 900 4307
rect 1548 4255 1554 4307
rect 894 4135 1554 4255
rect 894 4083 900 4135
rect 1548 4083 1554 4135
rect 894 3963 1554 4083
rect 894 3911 900 3963
rect 1548 3911 1554 3963
rect 894 3791 1554 3911
rect 894 3739 900 3791
rect 1548 3739 1554 3791
rect 894 3619 1554 3739
rect 894 3567 900 3619
rect 1548 3567 1554 3619
rect 894 3447 1554 3567
rect 894 3395 900 3447
rect 1548 3395 1554 3447
rect 894 3275 1554 3395
rect 894 3223 900 3275
rect 1548 3223 1554 3275
rect 894 3103 1554 3223
rect 894 3051 900 3103
rect 1548 3051 1554 3103
rect 894 2931 1554 3051
rect 894 2879 900 2931
rect 1548 2879 1554 2931
rect 894 2759 1554 2879
rect 894 2707 900 2759
rect 1548 2707 1554 2759
rect 894 2587 1554 2707
rect 894 2535 900 2587
rect 1548 2535 1554 2587
rect 894 2415 1554 2535
rect 894 2363 900 2415
rect 1548 2363 1554 2415
rect 894 2243 1554 2363
rect 894 2191 900 2243
rect 1548 2191 1554 2243
rect 894 2071 1554 2191
rect 894 2019 900 2071
rect 1548 2019 1554 2071
rect 894 1899 1554 2019
rect 894 1847 900 1899
rect 1548 1847 1554 1899
rect 894 1727 1554 1847
rect 894 1675 900 1727
rect 1548 1675 1554 1727
rect 894 1555 1554 1675
rect 894 1503 900 1555
rect 1548 1503 1554 1555
rect 894 1383 1554 1503
rect 894 1331 900 1383
rect 1548 1331 1554 1383
rect 894 1211 1554 1331
rect 894 1159 900 1211
rect 1548 1159 1554 1211
rect 894 1039 1554 1159
rect 894 987 900 1039
rect 1548 987 1554 1039
rect 894 867 1554 987
rect 894 815 900 867
rect 1548 815 1554 867
rect 894 695 1554 815
rect 894 643 900 695
rect 1548 643 1554 695
rect 894 523 1554 643
rect 894 471 900 523
rect 1548 471 1554 523
rect 894 351 1554 471
rect 894 299 900 351
rect 1548 299 1554 351
rect 894 179 1554 299
rect 894 127 900 179
rect 1548 127 1554 179
rect 1618 100069 1672 100075
rect 1618 163 1672 169
<< end >>
