VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_asw_1v8
  CLASS BLOCK ;
  FOREIGN tt_asw_1v8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 18.400 BY 21.760 ;
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.600 0.000 1.800 21.760 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 16.600 0.000 17.800 21.760 ;
    END
  END VPWR
  PIN mod
    DIRECTION INOUT ;
    USE ANALOG ;
    ANTENNADIFFAREA 5.675000 ;
    PORT
      LAYER met4 ;
        RECT 8.750 19.760 9.650 21.760 ;
    END
  END mod
  PIN bus
    DIRECTION INOUT ;
    USE ANALOG ;
    ANTENNADIFFAREA 5.675000 ;
    PORT
      LAYER met4 ;
        RECT 8.750 11.760 9.650 13.760 ;
    END
  END bus
  PIN ctrl
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.125000 ;
    PORT
      LAYER met3 ;
        RECT 4.450 20.860 4.750 21.760 ;
    END
  END ctrl
  OBS
      LAYER pwell ;
        RECT 2.500 15.000 4.610 19.600 ;
        RECT 4.850 17.250 5.300 17.550 ;
      LAYER nwell ;
        RECT 5.500 15.000 8.130 19.690 ;
        RECT 10.500 15.500 16.010 20.190 ;
      LAYER pwell ;
        RECT 2.500 8.000 4.610 12.600 ;
      LAYER nwell ;
        RECT 5.500 8.000 8.130 12.690 ;
      LAYER pwell ;
        RECT 10.500 9.700 14.090 14.300 ;
      LAYER li1 ;
        RECT 2.300 20.420 3.200 21.580 ;
        RECT 10.680 19.840 15.830 20.010 ;
        RECT 2.680 19.250 4.430 19.420 ;
        RECT 2.680 15.350 2.850 19.250 ;
        RECT 3.390 18.740 3.720 18.910 ;
        RECT 3.250 16.030 3.420 18.570 ;
        RECT 3.690 16.030 3.860 18.570 ;
        RECT 3.390 15.690 3.720 15.860 ;
        RECT 4.260 15.350 4.430 19.250 ;
        RECT 2.680 15.180 4.430 15.350 ;
        RECT 5.680 19.340 7.950 19.510 ;
        RECT 5.680 15.350 5.850 19.340 ;
        RECT 6.890 18.830 7.220 19.000 ;
        RECT 6.250 16.075 6.420 18.615 ;
        RECT 6.730 16.075 6.900 18.615 ;
        RECT 7.210 16.075 7.380 18.615 ;
        RECT 7.780 17.020 7.950 19.340 ;
        RECT 7.730 16.780 7.970 17.020 ;
        RECT 6.410 15.690 6.740 15.860 ;
        RECT 7.780 15.350 7.950 16.780 ;
        RECT 10.680 15.850 10.850 19.840 ;
        RECT 11.890 19.330 12.220 19.500 ;
        RECT 12.850 19.330 13.180 19.500 ;
        RECT 13.810 19.330 14.140 19.500 ;
        RECT 14.770 19.330 15.100 19.500 ;
        RECT 11.250 16.575 11.420 19.115 ;
        RECT 11.730 16.575 11.900 19.115 ;
        RECT 12.210 16.575 12.380 19.115 ;
        RECT 12.690 16.575 12.860 19.115 ;
        RECT 13.170 16.575 13.340 19.115 ;
        RECT 13.650 16.575 13.820 19.115 ;
        RECT 14.130 16.575 14.300 19.115 ;
        RECT 14.610 16.575 14.780 19.115 ;
        RECT 15.090 16.575 15.260 19.115 ;
        RECT 11.410 16.190 11.740 16.360 ;
        RECT 12.370 16.190 12.700 16.360 ;
        RECT 13.330 16.190 13.660 16.360 ;
        RECT 14.290 16.190 14.620 16.360 ;
        RECT 14.180 15.850 14.420 15.870 ;
        RECT 15.660 15.850 15.830 19.840 ;
        RECT 10.680 15.680 15.830 15.850 ;
        RECT 14.180 15.630 14.420 15.680 ;
        RECT 5.680 15.180 7.950 15.350 ;
        RECT 10.680 13.950 13.910 14.120 ;
        RECT 2.680 12.250 4.430 12.420 ;
        RECT 2.680 8.350 2.850 12.250 ;
        RECT 3.390 11.740 3.720 11.910 ;
        RECT 3.250 9.030 3.420 11.570 ;
        RECT 3.690 9.030 3.860 11.570 ;
        RECT 3.390 8.690 3.720 8.860 ;
        RECT 4.260 8.350 4.430 12.250 ;
        RECT 2.680 8.180 4.430 8.350 ;
        RECT 5.680 12.340 7.950 12.510 ;
        RECT 5.680 8.350 5.850 12.340 ;
        RECT 6.890 11.830 7.220 12.000 ;
        RECT 6.250 9.075 6.420 11.615 ;
        RECT 6.730 9.075 6.900 11.615 ;
        RECT 7.210 9.075 7.380 11.615 ;
        RECT 7.780 11.020 7.950 12.340 ;
        RECT 7.730 10.780 7.970 11.020 ;
        RECT 6.410 8.690 6.740 8.860 ;
        RECT 7.780 8.350 7.950 10.780 ;
        RECT 10.680 10.050 10.850 13.950 ;
        RECT 11.890 13.440 12.220 13.610 ;
        RECT 12.850 13.440 13.180 13.610 ;
        RECT 11.250 10.730 11.420 13.270 ;
        RECT 11.730 10.730 11.900 13.270 ;
        RECT 12.210 10.730 12.380 13.270 ;
        RECT 12.690 10.730 12.860 13.270 ;
        RECT 13.170 10.730 13.340 13.270 ;
        RECT 11.410 10.390 11.740 10.560 ;
        RECT 12.370 10.390 12.700 10.560 ;
        RECT 13.740 10.050 13.910 13.950 ;
        RECT 10.680 9.880 13.910 10.050 ;
        RECT 5.680 8.180 7.950 8.350 ;
      LAYER mcon ;
        RECT 2.400 20.700 3.100 21.300 ;
        RECT 3.470 18.740 3.640 18.910 ;
        RECT 3.250 16.110 3.420 18.490 ;
        RECT 3.690 16.110 3.860 18.490 ;
        RECT 3.470 15.690 3.640 15.860 ;
        RECT 6.970 18.830 7.140 19.000 ;
        RECT 6.250 16.155 6.420 18.535 ;
        RECT 6.730 16.155 6.900 18.535 ;
        RECT 7.210 16.155 7.380 18.535 ;
        RECT 7.730 16.780 7.970 17.020 ;
        RECT 6.490 15.690 6.660 15.860 ;
        RECT 11.970 19.330 12.140 19.500 ;
        RECT 12.930 19.330 13.100 19.500 ;
        RECT 13.890 19.330 14.060 19.500 ;
        RECT 14.850 19.330 15.020 19.500 ;
        RECT 11.250 16.655 11.420 19.035 ;
        RECT 11.730 16.655 11.900 19.035 ;
        RECT 12.210 16.655 12.380 19.035 ;
        RECT 12.690 16.655 12.860 19.035 ;
        RECT 13.170 16.655 13.340 19.035 ;
        RECT 13.650 16.655 13.820 19.035 ;
        RECT 14.130 16.655 14.300 19.035 ;
        RECT 14.610 16.655 14.780 19.035 ;
        RECT 15.090 16.655 15.260 19.035 ;
        RECT 11.490 16.190 11.660 16.360 ;
        RECT 12.450 16.190 12.620 16.360 ;
        RECT 13.410 16.190 13.580 16.360 ;
        RECT 14.370 16.190 14.540 16.360 ;
        RECT 3.470 11.740 3.640 11.910 ;
        RECT 3.250 9.110 3.420 11.490 ;
        RECT 3.690 9.110 3.860 11.490 ;
        RECT 3.470 8.690 3.640 8.860 ;
        RECT 6.970 11.830 7.140 12.000 ;
        RECT 6.250 9.155 6.420 11.535 ;
        RECT 6.730 9.155 6.900 11.535 ;
        RECT 7.210 9.155 7.380 11.535 ;
        RECT 7.730 10.780 7.970 11.020 ;
        RECT 6.490 8.690 6.660 8.860 ;
        RECT 11.970 13.440 12.140 13.610 ;
        RECT 12.930 13.440 13.100 13.610 ;
        RECT 11.250 10.810 11.420 13.190 ;
        RECT 11.730 10.810 11.900 13.190 ;
        RECT 12.210 10.810 12.380 13.190 ;
        RECT 12.690 10.810 12.860 13.190 ;
        RECT 13.170 10.810 13.340 13.190 ;
        RECT 11.490 10.390 11.660 10.560 ;
        RECT 12.450 10.390 12.620 10.560 ;
      LAYER met1 ;
        RECT 2.200 21.350 3.200 21.400 ;
        RECT 1.525 20.655 3.200 21.350 ;
        RECT 2.200 20.600 3.200 20.655 ;
        RECT 11.270 20.650 16.450 21.050 ;
        RECT 3.420 19.850 3.780 20.150 ;
        RECT 3.450 19.575 7.200 19.850 ;
        RECT 8.340 19.575 8.660 19.580 ;
        RECT 3.450 19.550 8.660 19.575 ;
        RECT 3.450 18.940 3.750 19.550 ;
        RECT 6.875 19.325 8.660 19.550 ;
        RECT 3.410 18.710 3.750 18.940 ;
        RECT 6.900 18.750 7.200 19.325 ;
        RECT 8.340 19.320 8.660 19.325 ;
        RECT 9.400 19.300 15.200 19.600 ;
        RECT 3.450 18.700 3.750 18.710 ;
        RECT 3.220 17.550 3.450 18.550 ;
        RECT 3.660 17.550 3.890 18.550 ;
        RECT 5.120 17.550 5.420 18.010 ;
        RECT 6.220 17.970 6.450 18.595 ;
        RECT 6.150 17.680 6.540 17.970 ;
        RECT 2.075 17.255 3.450 17.550 ;
        RECT 3.220 16.050 3.450 17.255 ;
        RECT 3.650 17.250 5.420 17.550 ;
        RECT 3.660 16.050 3.890 17.250 ;
        RECT 3.400 14.850 3.700 15.900 ;
        RECT 3.370 14.550 3.730 14.850 ;
        RECT 4.850 14.700 5.150 17.250 ;
        RECT 6.220 16.095 6.450 17.680 ;
        RECT 6.700 17.380 6.930 18.595 ;
        RECT 7.180 17.970 7.410 18.595 ;
        RECT 7.110 17.680 7.500 17.970 ;
        RECT 6.630 17.090 7.020 17.380 ;
        RECT 6.700 16.095 6.930 17.090 ;
        RECT 7.180 16.095 7.410 17.680 ;
        RECT 7.750 17.250 9.230 17.550 ;
        RECT 8.550 17.050 8.850 17.250 ;
        RECT 7.670 16.750 8.850 17.050 ;
        RECT 8.370 15.900 8.630 15.935 ;
        RECT 6.400 15.650 8.630 15.900 ;
        RECT 8.370 15.615 8.630 15.650 ;
        RECT 9.400 14.700 9.700 19.300 ;
        RECT 11.220 18.730 11.450 19.095 ;
        RECT 11.130 18.450 11.530 18.730 ;
        RECT 11.220 16.595 11.450 18.450 ;
        RECT 11.700 17.740 11.930 19.095 ;
        RECT 12.180 18.740 12.410 19.095 ;
        RECT 12.090 18.460 12.490 18.740 ;
        RECT 11.620 17.460 12.020 17.740 ;
        RECT 11.700 16.595 11.930 17.460 ;
        RECT 12.180 16.595 12.410 18.460 ;
        RECT 12.660 17.750 12.890 19.095 ;
        RECT 13.140 18.740 13.370 19.095 ;
        RECT 13.050 18.460 13.450 18.740 ;
        RECT 12.560 17.470 12.960 17.750 ;
        RECT 12.660 16.595 12.890 17.470 ;
        RECT 13.140 16.595 13.370 18.460 ;
        RECT 13.620 17.740 13.850 19.095 ;
        RECT 14.100 18.720 14.330 19.095 ;
        RECT 14.030 18.440 14.430 18.720 ;
        RECT 13.550 17.460 13.950 17.740 ;
        RECT 13.620 16.595 13.850 17.460 ;
        RECT 14.100 16.595 14.330 18.440 ;
        RECT 14.580 17.720 14.810 19.095 ;
        RECT 15.060 18.740 15.290 19.095 ;
        RECT 14.980 18.460 15.380 18.740 ;
        RECT 14.490 17.440 14.890 17.720 ;
        RECT 14.580 16.595 14.810 17.440 ;
        RECT 15.060 16.595 15.290 18.460 ;
        RECT 16.050 17.800 16.450 20.650 ;
        RECT 15.570 17.400 16.450 17.800 ;
        RECT 11.400 16.100 14.700 16.400 ;
        RECT 11.900 14.700 12.200 16.100 ;
        RECT 14.150 15.200 14.450 15.930 ;
        RECT 14.850 15.200 15.150 15.230 ;
        RECT 14.150 14.900 15.150 15.200 ;
        RECT 14.850 14.870 15.150 14.900 ;
        RECT 4.850 14.400 12.200 14.700 ;
        RECT 2.690 13.475 3.010 13.480 ;
        RECT 2.690 13.450 3.975 13.475 ;
        RECT 4.850 13.450 5.150 14.400 ;
        RECT 8.250 13.450 8.550 13.480 ;
        RECT 11.900 13.450 14.400 13.750 ;
        RECT 2.690 13.225 8.550 13.450 ;
        RECT 11.910 13.410 12.200 13.450 ;
        RECT 12.870 13.410 13.160 13.450 ;
        RECT 2.690 13.220 3.010 13.225 ;
        RECT 3.450 13.150 8.550 13.225 ;
        RECT 1.900 10.450 2.200 12.830 ;
        RECT 3.450 11.940 3.700 13.150 ;
        RECT 6.950 12.030 7.200 13.150 ;
        RECT 8.250 13.120 8.550 13.150 ;
        RECT 3.410 11.710 3.700 11.940 ;
        RECT 6.910 11.800 7.200 12.030 ;
        RECT 3.450 11.700 3.700 11.710 ;
        RECT 3.220 10.450 3.450 11.550 ;
        RECT 3.660 10.450 3.890 11.550 ;
        RECT 1.900 10.150 3.450 10.450 ;
        RECT 3.650 10.150 5.640 10.450 ;
        RECT 6.220 10.420 6.450 11.595 ;
        RECT 6.170 10.160 6.530 10.420 ;
        RECT 3.220 9.050 3.450 10.150 ;
        RECT 3.660 9.050 3.890 10.150 ;
        RECT 4.850 9.500 5.150 10.150 ;
        RECT 4.820 9.200 5.180 9.500 ;
        RECT 6.220 9.095 6.450 10.160 ;
        RECT 6.700 9.730 6.930 11.595 ;
        RECT 7.180 10.430 7.410 11.595 ;
        RECT 11.220 11.490 11.450 13.250 ;
        RECT 11.700 12.260 11.930 13.250 ;
        RECT 11.630 11.990 11.990 12.260 ;
        RECT 11.160 11.220 11.520 11.490 ;
        RECT 7.670 10.750 9.000 11.050 ;
        RECT 11.220 10.750 11.450 11.220 ;
        RECT 11.700 10.750 11.930 11.990 ;
        RECT 12.180 11.490 12.410 13.250 ;
        RECT 12.660 12.260 12.890 13.250 ;
        RECT 12.600 11.990 12.960 12.260 ;
        RECT 12.110 11.220 12.470 11.490 ;
        RECT 12.180 10.750 12.410 11.220 ;
        RECT 12.660 10.750 12.890 11.990 ;
        RECT 13.140 11.480 13.370 13.250 ;
        RECT 13.090 11.210 13.450 11.480 ;
        RECT 13.140 10.750 13.370 11.210 ;
        RECT 8.700 10.450 9.000 10.750 ;
        RECT 7.130 10.170 7.490 10.430 ;
        RECT 6.630 9.470 6.990 9.730 ;
        RECT 6.700 9.095 6.930 9.470 ;
        RECT 7.180 9.095 7.410 10.170 ;
        RECT 8.200 10.150 9.000 10.450 ;
        RECT 11.400 10.300 12.700 10.600 ;
        RECT 8.200 9.750 8.500 10.150 ;
        RECT 7.700 9.450 8.500 9.750 ;
        RECT 8.700 8.950 9.000 10.150 ;
        RECT 11.900 9.270 12.200 10.300 ;
        RECT 13.000 9.600 13.300 9.630 ;
        RECT 14.100 9.600 14.400 13.450 ;
        RECT 13.000 9.300 14.400 9.600 ;
        RECT 13.000 9.270 13.300 9.300 ;
        RECT 14.750 8.950 15.050 13.080 ;
        RECT 16.050 11.550 16.450 17.400 ;
        RECT 15.320 11.150 16.450 11.550 ;
        RECT 3.450 8.890 3.700 8.900 ;
        RECT 3.410 8.660 3.700 8.890 ;
        RECT 2.690 7.875 3.010 7.880 ;
        RECT 3.450 7.875 3.700 8.660 ;
        RECT 2.690 7.625 3.700 7.875 ;
        RECT 2.690 7.620 3.010 7.625 ;
        RECT 3.450 7.600 3.700 7.625 ;
        RECT 6.400 8.890 6.700 8.900 ;
        RECT 6.400 8.660 6.720 8.890 ;
        RECT 6.400 7.100 6.700 8.660 ;
        RECT 8.700 8.650 15.100 8.950 ;
        RECT 8.250 7.100 8.550 8.380 ;
        RECT 6.400 6.800 8.550 7.100 ;
      LAYER via ;
        RECT 1.555 20.655 2.250 21.350 ;
        RECT 11.300 20.650 11.700 21.050 ;
        RECT 3.450 19.850 3.750 20.150 ;
        RECT 8.370 19.320 8.630 19.580 ;
        RECT 5.120 17.680 5.420 17.980 ;
        RECT 6.200 17.680 6.490 17.970 ;
        RECT 2.105 17.255 2.400 17.550 ;
        RECT 3.400 14.550 3.700 14.850 ;
        RECT 7.160 17.680 7.450 17.970 ;
        RECT 6.680 17.090 6.970 17.380 ;
        RECT 7.780 17.250 8.080 17.550 ;
        RECT 8.900 17.250 9.200 17.550 ;
        RECT 8.370 15.645 8.630 15.905 ;
        RECT 11.180 18.450 11.480 18.730 ;
        RECT 12.140 18.460 12.440 18.740 ;
        RECT 11.670 17.460 11.970 17.740 ;
        RECT 13.100 18.460 13.400 18.740 ;
        RECT 12.610 17.470 12.910 17.750 ;
        RECT 14.080 18.440 14.380 18.720 ;
        RECT 13.600 17.460 13.900 17.740 ;
        RECT 15.030 18.460 15.330 18.740 ;
        RECT 14.540 17.440 14.840 17.720 ;
        RECT 15.600 17.400 16.000 17.800 ;
        RECT 14.850 14.900 15.150 15.200 ;
        RECT 2.720 13.220 2.980 13.480 ;
        RECT 8.250 13.150 8.550 13.450 ;
        RECT 1.900 12.500 2.200 12.800 ;
        RECT 5.310 10.150 5.610 10.450 ;
        RECT 6.220 10.160 6.480 10.420 ;
        RECT 4.850 9.200 5.150 9.500 ;
        RECT 11.680 11.990 11.940 12.260 ;
        RECT 11.210 11.220 11.470 11.490 ;
        RECT 12.650 11.990 12.910 12.260 ;
        RECT 12.160 11.220 12.420 11.490 ;
        RECT 13.140 11.210 13.400 11.480 ;
        RECT 7.180 10.170 7.440 10.430 ;
        RECT 6.680 9.470 6.940 9.730 ;
        RECT 7.730 9.450 8.030 9.750 ;
        RECT 11.900 9.300 12.200 9.600 ;
        RECT 14.750 12.750 15.050 13.050 ;
        RECT 15.350 11.150 15.750 11.550 ;
        RECT 2.720 7.620 2.980 7.880 ;
        RECT 8.250 8.050 8.550 8.350 ;
      LAYER met2 ;
        RECT 1.555 21.350 2.250 21.380 ;
        RECT 1.010 20.655 2.250 21.350 ;
        RECT 11.300 21.050 11.700 21.080 ;
        RECT 1.555 20.625 2.250 20.655 ;
        RECT 3.450 20.150 3.750 20.745 ;
        RECT 10.055 20.650 11.700 21.050 ;
        RECT 11.300 20.620 11.700 20.650 ;
        RECT 3.450 19.850 4.650 20.150 ;
        RECT 3.450 19.820 3.750 19.850 ;
        RECT 1.360 17.550 1.750 17.555 ;
        RECT 2.105 17.550 2.400 17.580 ;
        RECT 1.360 17.255 2.400 17.550 ;
        RECT 2.105 17.225 2.400 17.255 ;
        RECT 3.400 14.850 3.700 14.880 ;
        RECT 4.350 14.850 4.650 19.850 ;
        RECT 8.370 19.290 8.630 19.610 ;
        RECT 6.200 17.980 6.490 18.020 ;
        RECT 7.160 17.980 7.450 18.020 ;
        RECT 5.090 17.680 7.600 17.980 ;
        RECT 6.200 17.630 6.490 17.680 ;
        RECT 7.160 17.630 7.450 17.680 ;
        RECT 6.680 17.390 6.970 17.430 ;
        RECT 7.780 17.390 8.080 17.580 ;
        RECT 6.060 17.090 8.080 17.390 ;
        RECT 6.680 17.040 6.970 17.090 ;
        RECT 8.375 15.905 8.625 19.290 ;
        RECT 11.180 18.775 11.480 18.780 ;
        RECT 12.140 18.775 12.440 18.790 ;
        RECT 13.100 18.775 13.400 18.790 ;
        RECT 15.030 18.775 15.330 18.790 ;
        RECT 10.075 18.425 15.425 18.775 ;
        RECT 8.900 17.550 9.200 17.580 ;
        RECT 8.900 17.250 9.745 17.550 ;
        RECT 8.900 17.220 9.200 17.250 ;
        RECT 8.340 15.645 8.660 15.905 ;
        RECT 3.400 14.550 4.650 14.850 ;
        RECT 3.400 14.520 3.700 14.550 ;
        RECT 2.720 13.190 2.980 13.510 ;
        RECT 1.055 12.500 2.230 12.800 ;
        RECT 2.725 7.910 2.975 13.190 ;
        RECT 8.220 13.150 8.580 13.450 ;
        RECT 5.310 10.450 5.610 10.480 ;
        RECT 6.220 10.450 6.480 10.470 ;
        RECT 7.180 10.450 7.440 10.480 ;
        RECT 5.310 10.150 7.510 10.450 ;
        RECT 5.310 10.120 5.610 10.150 ;
        RECT 6.220 10.110 6.480 10.150 ;
        RECT 7.180 10.120 7.440 10.150 ;
        RECT 6.680 9.750 6.940 9.780 ;
        RECT 7.730 9.750 8.030 9.780 ;
        RECT 2.720 7.590 2.980 7.910 ;
        RECT 4.850 7.800 5.150 9.530 ;
        RECT 6.060 9.450 8.030 9.750 ;
        RECT 6.680 9.420 6.940 9.450 ;
        RECT 7.730 9.420 8.030 9.450 ;
        RECT 8.250 8.350 8.550 13.150 ;
        RECT 10.075 13.075 10.425 18.425 ;
        RECT 11.180 18.400 11.480 18.425 ;
        RECT 12.140 18.410 12.440 18.425 ;
        RECT 13.100 18.410 13.400 18.425 ;
        RECT 14.080 18.390 14.380 18.425 ;
        RECT 15.030 18.410 15.330 18.425 ;
        RECT 15.600 17.800 16.000 17.830 ;
        RECT 11.100 17.400 16.000 17.800 ;
        RECT 14.540 17.390 14.840 17.400 ;
        RECT 15.600 17.370 16.000 17.400 ;
        RECT 15.610 15.200 15.890 15.235 ;
        RECT 14.820 14.900 15.900 15.200 ;
        RECT 15.610 14.865 15.890 14.900 ;
        RECT 10.030 12.725 10.470 13.075 ;
        RECT 14.720 12.750 15.895 13.050 ;
        RECT 10.075 12.300 10.425 12.725 ;
        RECT 11.680 12.300 11.940 12.310 ;
        RECT 12.650 12.300 12.910 12.310 ;
        RECT 10.045 11.950 13.375 12.300 ;
        RECT 11.680 11.940 11.940 11.950 ;
        RECT 12.650 11.940 12.910 11.950 ;
        RECT 15.350 11.550 15.750 11.580 ;
        RECT 10.700 11.150 15.750 11.550 ;
        RECT 15.350 11.120 15.750 11.150 ;
        RECT 11.870 9.300 13.330 9.600 ;
        RECT 8.220 8.050 8.580 8.350 ;
        RECT 11.900 7.800 12.200 9.300 ;
        RECT 4.850 7.500 12.200 7.800 ;
      LAYER via2 ;
        RECT 1.055 20.655 1.750 21.350 ;
        RECT 3.450 20.400 3.750 20.700 ;
        RECT 10.100 20.650 10.500 21.050 ;
        RECT 1.405 17.255 1.705 17.555 ;
        RECT 9.400 17.250 9.700 17.550 ;
        RECT 1.100 12.500 1.400 12.800 ;
        RECT 15.610 14.910 15.890 15.190 ;
        RECT 10.075 12.725 10.425 13.075 ;
        RECT 15.550 12.750 15.850 13.050 ;
      LAYER met3 ;
        RECT 0.600 11.760 1.800 21.760 ;
        RECT 3.450 21.200 4.450 21.500 ;
        RECT 3.450 20.725 3.750 21.200 ;
        RECT 8.750 21.050 9.650 21.760 ;
        RECT 10.075 21.050 10.525 21.075 ;
        RECT 3.425 20.375 3.775 20.725 ;
        RECT 4.450 20.650 4.750 20.860 ;
        RECT 8.750 20.650 10.525 21.050 ;
        RECT 8.750 19.760 9.650 20.650 ;
        RECT 10.075 20.625 10.525 20.650 ;
        RECT 9.375 17.550 9.725 17.575 ;
        RECT 16.600 17.550 17.800 21.760 ;
        RECT 9.375 17.250 17.800 17.550 ;
        RECT 9.375 17.225 9.725 17.250 ;
        RECT 15.585 15.200 15.915 15.215 ;
        RECT 16.600 15.200 17.800 17.250 ;
        RECT 15.585 14.900 17.800 15.200 ;
        RECT 15.585 14.885 15.915 14.900 ;
        RECT 8.750 13.075 9.650 13.760 ;
        RECT 15.540 13.510 15.860 13.890 ;
        RECT 10.050 13.075 10.450 13.100 ;
        RECT 15.550 13.075 15.850 13.510 ;
        RECT 8.750 12.725 10.450 13.075 ;
        RECT 15.525 12.725 15.875 13.075 ;
        RECT 8.750 11.760 9.650 12.725 ;
        RECT 10.050 12.700 10.450 12.725 ;
        RECT 16.600 11.760 17.800 14.900 ;
      LAYER via3 ;
        RECT 0.630 11.790 1.770 21.730 ;
        RECT 8.780 19.790 9.620 21.730 ;
        RECT 8.780 11.790 9.620 13.730 ;
        RECT 15.540 13.540 15.860 13.860 ;
        RECT 16.630 11.790 17.770 21.730 ;
      LAYER met4 ;
        RECT 15.535 13.850 15.865 13.865 ;
        RECT 15.535 13.550 16.600 13.850 ;
        RECT 15.535 13.535 15.865 13.550 ;
  END
END tt_asw_1v8
END LIBRARY

