magic
tech sky130A
magscale 1 2
timestamp 1718383489
<< metal2 >>
rect 299 1115 1379 1120
rect 299 5 308 1115
rect 1370 5 1379 1115
rect 299 0 1379 5
rect 1459 1115 2539 1120
rect 1459 5 1633 1115
rect 2530 5 2539 1115
rect 1459 0 2539 5
<< via2 >>
rect 308 5 1370 1115
rect 1633 5 2530 1115
<< metal3 >>
rect 299 1119 1504 1120
rect 299 1115 686 1119
rect 299 5 308 1115
rect 299 1 686 5
rect 1498 1 1504 1119
rect 299 0 1504 1
rect 1624 1119 2760 1120
rect 1624 1115 1776 1119
rect 1624 5 1633 1115
rect 1624 1 1776 5
rect 2754 1 2760 1119
rect 1624 0 2760 1
<< via3 >>
rect 686 1115 1498 1119
rect 686 5 1370 1115
rect 1370 5 1498 1115
rect 686 1 1498 5
rect 1776 1115 2754 1119
rect 1776 5 2530 1115
rect 2530 5 2754 1115
rect 1776 1 2754 5
<< metal4 >>
rect 0 0 240 1120
rect 340 0 580 1120
rect 680 1119 1670 1120
rect 680 1 686 1119
rect 1498 1 1670 1119
rect 680 0 1670 1
rect 1770 1119 2760 1120
rect 1770 1 1776 1119
rect 2754 1 2760 1119
rect 1770 0 2760 1
<< end >>
