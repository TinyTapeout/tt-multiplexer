magic
tech sky130A
magscale 1 2
timestamp 1712317355
<< nwell >>
rect -263 -369 263 369
<< pmos >>
rect -63 -150 -33 150
rect 33 -150 63 150
<< pdiff >>
rect -125 138 -63 150
rect -125 -138 -113 138
rect -79 -138 -63 138
rect -125 -150 -63 -138
rect -33 138 33 150
rect -33 -138 -17 138
rect 17 -138 33 138
rect -33 -150 33 -138
rect 63 138 125 150
rect 63 -138 79 138
rect 113 -138 125 138
rect 63 -150 125 -138
<< pdiffc >>
rect -113 -138 -79 138
rect -17 -138 17 138
rect 79 -138 113 138
<< nsubdiff >>
rect -227 299 -131 333
rect 131 299 227 333
rect -227 237 -193 299
rect 193 237 227 299
rect -227 -299 -193 -237
rect 193 -299 227 -237
rect -227 -333 -131 -299
rect 131 -333 227 -299
<< nsubdiffcont >>
rect -131 299 131 333
rect -227 -237 -193 237
rect 193 -237 227 237
rect -131 -333 131 -299
<< poly >>
rect -82 231 82 248
rect -82 197 -65 231
rect -31 197 31 231
rect 65 197 82 231
rect -82 180 82 197
rect -63 150 -33 180
rect 33 150 63 180
rect -63 -180 -33 -150
rect 33 -180 63 -150
rect -82 -197 82 -180
rect -82 -231 -65 -197
rect -31 -231 31 -197
rect 65 -231 82 -197
rect -82 -248 82 -231
<< polycont >>
rect -65 197 -31 231
rect 31 197 65 231
rect -65 -231 -31 -197
rect 31 -231 65 -197
<< locali >>
rect -227 299 -131 333
rect 131 299 227 333
rect -227 237 -193 299
rect 193 237 227 299
rect -82 231 82 232
rect -82 197 -65 231
rect -31 197 31 231
rect 65 197 82 231
rect -82 196 82 197
rect -113 138 -79 154
rect -113 -154 -79 -138
rect -17 138 17 154
rect -17 -154 17 -138
rect 79 138 113 154
rect 79 -154 113 -138
rect -82 -197 82 -196
rect -82 -231 -65 -197
rect -31 -231 31 -197
rect 65 -231 82 -197
rect -82 -232 82 -231
rect -227 -299 -193 -237
rect 193 -299 227 -237
rect -227 -333 -131 -299
rect 131 -333 227 -299
<< viali >>
rect -65 197 -31 231
rect 31 197 65 231
rect -113 -138 -79 138
rect -17 -138 17 138
rect 79 -138 113 138
rect -65 -231 -31 -197
rect 31 -231 65 -197
<< metal1 >>
rect -82 231 82 238
rect -82 197 -65 231
rect -31 197 31 231
rect 65 197 82 231
rect -82 190 82 197
rect -119 138 -73 150
rect -119 -138 -113 138
rect -79 -138 -73 138
rect -119 -150 -73 -138
rect -23 138 23 150
rect -23 -138 -17 138
rect 17 -138 23 138
rect -23 -150 23 -138
rect 73 138 119 150
rect 73 -138 79 138
rect 113 -138 119 138
rect 73 -150 119 -138
rect -82 -197 82 -190
rect -82 -231 -65 -197
rect -31 -231 82 -197
rect -82 -238 82 -231
<< properties >>
string FIXED_BBOX -210 -316 210 316
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.5 l 0.15 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
