magic
tech sky130A
magscale 1 2
timestamp 1712480545
<< error_p >>
rect -415 522 -353 528
rect -287 522 -225 528
rect -159 522 -97 528
rect -31 522 31 528
rect 97 522 159 528
rect 225 522 287 528
rect 353 522 415 528
rect -415 488 -403 522
rect -287 488 -275 522
rect -159 488 -147 522
rect -31 488 -19 522
rect 97 488 109 522
rect 225 488 237 522
rect 353 488 365 522
rect -415 482 -353 488
rect -287 482 -225 488
rect -159 482 -97 488
rect -31 482 31 488
rect 97 482 159 488
rect 225 482 287 488
rect 353 482 415 488
rect -415 -488 -353 -482
rect -287 -488 -225 -482
rect -159 -488 -97 -482
rect -31 -488 31 -482
rect 97 -488 159 -482
rect 225 -488 287 -482
rect 353 -488 415 -482
rect -415 -522 -403 -488
rect -287 -522 -275 -488
rect -159 -522 -147 -488
rect -31 -522 -19 -488
rect 97 -522 109 -488
rect 225 -522 237 -488
rect 353 -522 365 -488
rect -415 -528 -353 -522
rect -287 -528 -225 -522
rect -159 -528 -97 -522
rect -31 -528 31 -522
rect 97 -528 159 -522
rect 225 -528 287 -522
rect 353 -528 415 -522
<< pwell >>
rect -615 -660 615 660
<< nmoslvt >>
rect -419 -450 -349 450
rect -291 -450 -221 450
rect -163 -450 -93 450
rect -35 -450 35 450
rect 93 -450 163 450
rect 221 -450 291 450
rect 349 -450 419 450
<< ndiff >>
rect -477 438 -419 450
rect -477 -438 -465 438
rect -431 -438 -419 438
rect -477 -450 -419 -438
rect -349 438 -291 450
rect -349 -438 -337 438
rect -303 -438 -291 438
rect -349 -450 -291 -438
rect -221 438 -163 450
rect -221 -438 -209 438
rect -175 -438 -163 438
rect -221 -450 -163 -438
rect -93 438 -35 450
rect -93 -438 -81 438
rect -47 -438 -35 438
rect -93 -450 -35 -438
rect 35 438 93 450
rect 35 -438 47 438
rect 81 -438 93 438
rect 35 -450 93 -438
rect 163 438 221 450
rect 163 -438 175 438
rect 209 -438 221 438
rect 163 -450 221 -438
rect 291 438 349 450
rect 291 -438 303 438
rect 337 -438 349 438
rect 291 -450 349 -438
rect 419 438 477 450
rect 419 -438 431 438
rect 465 -438 477 438
rect 419 -450 477 -438
<< ndiffc >>
rect -465 -438 -431 438
rect -337 -438 -303 438
rect -209 -438 -175 438
rect -81 -438 -47 438
rect 47 -438 81 438
rect 175 -438 209 438
rect 303 -438 337 438
rect 431 -438 465 438
<< psubdiff >>
rect -579 590 -483 624
rect 483 590 579 624
rect -579 528 -545 590
rect 545 528 579 590
rect -579 -590 -545 -528
rect 545 -590 579 -528
rect -579 -624 -483 -590
rect 483 -624 579 -590
<< psubdiffcont >>
rect -483 590 483 624
rect -579 -528 -545 528
rect 545 -528 579 528
rect -483 -624 483 -590
<< poly >>
rect -419 522 -349 538
rect -419 488 -403 522
rect -365 488 -349 522
rect -419 450 -349 488
rect -291 522 -221 538
rect -291 488 -275 522
rect -237 488 -221 522
rect -291 450 -221 488
rect -163 522 -93 538
rect -163 488 -147 522
rect -109 488 -93 522
rect -163 450 -93 488
rect -35 522 35 538
rect -35 488 -19 522
rect 19 488 35 522
rect -35 450 35 488
rect 93 522 163 538
rect 93 488 109 522
rect 147 488 163 522
rect 93 450 163 488
rect 221 522 291 538
rect 221 488 237 522
rect 275 488 291 522
rect 221 450 291 488
rect 349 522 419 538
rect 349 488 365 522
rect 403 488 419 522
rect 349 450 419 488
rect -419 -488 -349 -450
rect -419 -522 -403 -488
rect -365 -522 -349 -488
rect -419 -538 -349 -522
rect -291 -488 -221 -450
rect -291 -522 -275 -488
rect -237 -522 -221 -488
rect -291 -538 -221 -522
rect -163 -488 -93 -450
rect -163 -522 -147 -488
rect -109 -522 -93 -488
rect -163 -538 -93 -522
rect -35 -488 35 -450
rect -35 -522 -19 -488
rect 19 -522 35 -488
rect -35 -538 35 -522
rect 93 -488 163 -450
rect 93 -522 109 -488
rect 147 -522 163 -488
rect 93 -538 163 -522
rect 221 -488 291 -450
rect 221 -522 237 -488
rect 275 -522 291 -488
rect 221 -538 291 -522
rect 349 -488 419 -450
rect 349 -522 365 -488
rect 403 -522 419 -488
rect 349 -538 419 -522
<< polycont >>
rect -403 488 -365 522
rect -275 488 -237 522
rect -147 488 -109 522
rect -19 488 19 522
rect 109 488 147 522
rect 237 488 275 522
rect 365 488 403 522
rect -403 -522 -365 -488
rect -275 -522 -237 -488
rect -147 -522 -109 -488
rect -19 -522 19 -488
rect 109 -522 147 -488
rect 237 -522 275 -488
rect 365 -522 403 -488
<< locali >>
rect -579 590 -483 624
rect 483 590 579 624
rect -579 528 -545 590
rect 545 528 579 590
rect -419 488 -403 522
rect -365 488 -349 522
rect -291 488 -275 522
rect -237 488 -221 522
rect -163 488 -147 522
rect -109 488 -93 522
rect -35 488 -19 522
rect 19 488 35 522
rect 93 488 109 522
rect 147 488 163 522
rect 221 488 237 522
rect 275 488 291 522
rect 349 488 365 522
rect 403 488 419 522
rect -465 438 -431 454
rect -465 -454 -431 -438
rect -337 438 -303 454
rect -337 -454 -303 -438
rect -209 438 -175 454
rect -209 -454 -175 -438
rect -81 438 -47 454
rect -81 -454 -47 -438
rect 47 438 81 454
rect 47 -454 81 -438
rect 175 438 209 454
rect 175 -454 209 -438
rect 303 438 337 454
rect 303 -454 337 -438
rect 431 438 465 454
rect 431 -454 465 -438
rect -419 -522 -403 -488
rect -365 -522 -349 -488
rect -291 -522 -275 -488
rect -237 -522 -221 -488
rect -163 -522 -147 -488
rect -109 -522 -93 -488
rect -35 -522 -19 -488
rect 19 -522 35 -488
rect 93 -522 109 -488
rect 147 -522 163 -488
rect 221 -522 237 -488
rect 275 -522 291 -488
rect 349 -522 365 -488
rect 403 -522 419 -488
rect -579 -590 -545 -528
rect 545 -590 579 -528
rect -579 -624 -483 -590
rect 483 -624 579 -590
<< viali >>
rect -403 488 -365 522
rect -275 488 -237 522
rect -147 488 -109 522
rect -19 488 19 522
rect 109 488 147 522
rect 237 488 275 522
rect 365 488 403 522
rect -465 -438 -431 438
rect -337 -438 -303 438
rect -209 -438 -175 438
rect -81 -438 -47 438
rect 47 -438 81 438
rect 175 -438 209 438
rect 303 -438 337 438
rect 431 -438 465 438
rect -403 -522 -365 -488
rect -275 -522 -237 -488
rect -147 -522 -109 -488
rect -19 -522 19 -488
rect 109 -522 147 -488
rect 237 -522 275 -488
rect 365 -522 403 -488
<< metal1 >>
rect -415 522 -353 528
rect -415 488 -403 522
rect -365 488 -353 522
rect -415 482 -353 488
rect -287 522 -225 528
rect -287 488 -275 522
rect -237 488 -225 522
rect -287 482 -225 488
rect -159 522 -97 528
rect -159 488 -147 522
rect -109 488 -97 522
rect -159 482 -97 488
rect -31 522 31 528
rect -31 488 -19 522
rect 19 488 31 522
rect -31 482 31 488
rect 97 522 159 528
rect 97 488 109 522
rect 147 488 159 522
rect 97 482 159 488
rect 225 522 287 528
rect 225 488 237 522
rect 275 488 287 522
rect 225 482 287 488
rect 353 522 415 528
rect 353 488 365 522
rect 403 488 415 522
rect 353 482 415 488
rect -471 438 -425 450
rect -471 -438 -465 438
rect -431 -438 -425 438
rect -471 -450 -425 -438
rect -343 438 -297 450
rect -343 -438 -337 438
rect -303 -438 -297 438
rect -343 -450 -297 -438
rect -215 438 -169 450
rect -215 -438 -209 438
rect -175 -438 -169 438
rect -215 -450 -169 -438
rect -87 438 -41 450
rect -87 -438 -81 438
rect -47 -438 -41 438
rect -87 -450 -41 -438
rect 41 438 87 450
rect 41 -438 47 438
rect 81 -438 87 438
rect 41 -450 87 -438
rect 169 438 215 450
rect 169 -438 175 438
rect 209 -438 215 438
rect 169 -450 215 -438
rect 297 438 343 450
rect 297 -438 303 438
rect 337 -438 343 438
rect 297 -450 343 -438
rect 425 438 471 450
rect 425 -438 431 438
rect 465 -438 471 438
rect 425 -450 471 -438
rect -415 -488 -353 -482
rect -415 -522 -403 -488
rect -365 -522 -353 -488
rect -415 -528 -353 -522
rect -287 -488 -225 -482
rect -287 -522 -275 -488
rect -237 -522 -225 -488
rect -287 -528 -225 -522
rect -159 -488 -97 -482
rect -159 -522 -147 -488
rect -109 -522 -97 -488
rect -159 -528 -97 -522
rect -31 -488 31 -482
rect -31 -522 -19 -488
rect 19 -522 31 -488
rect -31 -528 31 -522
rect 97 -488 159 -482
rect 97 -522 109 -488
rect 147 -522 159 -488
rect 97 -528 159 -522
rect 225 -488 287 -482
rect 225 -522 237 -488
rect 275 -522 287 -488
rect 225 -528 287 -522
rect 353 -488 415 -482
rect 353 -522 365 -488
rect 403 -522 415 -488
rect 353 -528 415 -522
<< properties >>
string FIXED_BBOX -562 -607 562 607
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 4.5 l 0.350 m 1 nf 7 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
