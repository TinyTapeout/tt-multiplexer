magic
tech sky130A
magscale 1 2
timestamp 1718382556
<< nwell >>
rect 0 0 2686 43110
<< mvpmos >>
rect 232 42799 2532 42899
rect 232 42643 2532 42743
rect 232 42487 2532 42587
rect 232 42331 2532 42431
rect 232 42175 2532 42275
rect 232 42019 2532 42119
rect 232 41863 2532 41963
rect 232 41707 2532 41807
rect 232 41551 2532 41651
rect 232 41395 2532 41495
rect 232 41239 2532 41339
rect 232 41083 2532 41183
rect 232 40927 2532 41027
rect 232 40771 2532 40871
rect 232 40615 2532 40715
rect 232 40459 2532 40559
rect 232 40303 2532 40403
rect 232 40147 2532 40247
rect 232 39991 2532 40091
rect 232 39835 2532 39935
rect 232 39679 2532 39779
rect 232 39523 2532 39623
rect 232 39367 2532 39467
rect 232 39211 2532 39311
rect 232 39055 2532 39155
rect 232 38899 2532 38999
rect 232 38743 2532 38843
rect 232 38587 2532 38687
rect 232 38431 2532 38531
rect 232 38275 2532 38375
rect 232 38119 2532 38219
rect 232 37963 2532 38063
rect 232 37807 2532 37907
rect 232 37651 2532 37751
rect 232 37495 2532 37595
rect 232 37339 2532 37439
rect 232 37183 2532 37283
rect 232 37027 2532 37127
rect 232 36871 2532 36971
rect 232 36715 2532 36815
rect 232 36559 2532 36659
rect 232 36403 2532 36503
rect 232 36247 2532 36347
rect 232 36091 2532 36191
rect 232 35935 2532 36035
rect 232 35779 2532 35879
rect 232 35623 2532 35723
rect 232 35467 2532 35567
rect 232 35311 2532 35411
rect 232 35155 2532 35255
rect 232 34999 2532 35099
rect 232 34843 2532 34943
rect 232 34687 2532 34787
rect 232 34531 2532 34631
rect 232 34375 2532 34475
rect 232 34219 2532 34319
rect 232 34063 2532 34163
rect 232 33907 2532 34007
rect 232 33751 2532 33851
rect 232 33595 2532 33695
rect 232 33439 2532 33539
rect 232 33283 2532 33383
rect 232 33127 2532 33227
rect 232 32971 2532 33071
rect 232 32815 2532 32915
rect 232 32659 2532 32759
rect 232 32503 2532 32603
rect 232 32347 2532 32447
rect 232 32191 2532 32291
rect 232 32035 2532 32135
rect 232 31879 2532 31979
rect 232 31723 2532 31823
rect 232 31567 2532 31667
rect 232 31411 2532 31511
rect 232 31255 2532 31355
rect 232 31099 2532 31199
rect 232 30943 2532 31043
rect 232 30787 2532 30887
rect 232 30631 2532 30731
rect 232 30475 2532 30575
rect 232 30319 2532 30419
rect 232 30163 2532 30263
rect 232 30007 2532 30107
rect 232 29851 2532 29951
rect 232 29695 2532 29795
rect 232 29539 2532 29639
rect 232 29383 2532 29483
rect 232 29227 2532 29327
rect 232 29071 2532 29171
rect 232 28915 2532 29015
rect 232 28759 2532 28859
rect 232 28603 2532 28703
rect 232 28447 2532 28547
rect 232 28291 2532 28391
rect 232 28135 2532 28235
rect 232 27979 2532 28079
rect 232 27823 2532 27923
rect 232 27667 2532 27767
rect 232 27511 2532 27611
rect 232 27355 2532 27455
rect 232 27199 2532 27299
rect 232 27043 2532 27143
rect 232 26887 2532 26987
rect 232 26731 2532 26831
rect 232 26575 2532 26675
rect 232 26419 2532 26519
rect 232 26263 2532 26363
rect 232 26107 2532 26207
rect 232 25951 2532 26051
rect 232 25795 2532 25895
rect 232 25639 2532 25739
rect 232 25483 2532 25583
rect 232 25327 2532 25427
rect 232 25171 2532 25271
rect 232 25015 2532 25115
rect 232 24859 2532 24959
rect 232 24703 2532 24803
rect 232 24547 2532 24647
rect 232 24391 2532 24491
rect 232 24235 2532 24335
rect 232 24079 2532 24179
rect 232 23923 2532 24023
rect 232 23767 2532 23867
rect 232 23611 2532 23711
rect 232 23455 2532 23555
rect 232 23299 2532 23399
rect 232 23143 2532 23243
rect 232 22987 2532 23087
rect 232 22831 2532 22931
rect 232 22675 2532 22775
rect 232 22519 2532 22619
rect 232 22363 2532 22463
rect 232 22207 2532 22307
rect 232 22051 2532 22151
rect 232 21895 2532 21995
rect 232 21739 2532 21839
rect 232 21583 2532 21683
rect 232 21427 2532 21527
rect 232 21271 2532 21371
rect 232 21115 2532 21215
rect 232 20959 2532 21059
rect 232 20803 2532 20903
rect 232 20647 2532 20747
rect 232 20491 2532 20591
rect 232 20335 2532 20435
rect 232 20179 2532 20279
rect 232 20023 2532 20123
rect 232 19867 2532 19967
rect 232 19711 2532 19811
rect 232 19555 2532 19655
rect 232 19399 2532 19499
rect 232 19243 2532 19343
rect 232 19087 2532 19187
rect 232 18931 2532 19031
rect 232 18775 2532 18875
rect 232 18619 2532 18719
rect 232 18463 2532 18563
rect 232 18307 2532 18407
rect 232 18151 2532 18251
rect 232 17995 2532 18095
rect 232 17839 2532 17939
rect 232 17683 2532 17783
rect 232 17527 2532 17627
rect 232 17371 2532 17471
rect 232 17215 2532 17315
rect 232 17059 2532 17159
rect 232 16903 2532 17003
rect 232 16747 2532 16847
rect 232 16591 2532 16691
rect 232 16435 2532 16535
rect 232 16279 2532 16379
rect 232 16123 2532 16223
rect 232 15967 2532 16067
rect 232 15811 2532 15911
rect 232 15655 2532 15755
rect 232 15499 2532 15599
rect 232 15343 2532 15443
rect 232 15187 2532 15287
rect 232 15031 2532 15131
rect 232 14875 2532 14975
rect 232 14719 2532 14819
rect 232 14563 2532 14663
rect 232 14407 2532 14507
rect 232 14251 2532 14351
rect 232 14095 2532 14195
rect 232 13939 2532 14039
rect 232 13783 2532 13883
rect 232 13627 2532 13727
rect 232 13471 2532 13571
rect 232 13315 2532 13415
rect 232 13159 2532 13259
rect 232 13003 2532 13103
rect 232 12847 2532 12947
rect 232 12691 2532 12791
rect 232 12535 2532 12635
rect 232 12379 2532 12479
rect 232 12223 2532 12323
rect 232 12067 2532 12167
rect 232 11911 2532 12011
rect 232 11755 2532 11855
rect 232 11599 2532 11699
rect 232 11443 2532 11543
rect 232 11287 2532 11387
rect 232 11131 2532 11231
rect 232 10975 2532 11075
rect 232 10819 2532 10919
rect 232 10663 2532 10763
rect 232 10507 2532 10607
rect 232 10351 2532 10451
rect 232 10195 2532 10295
rect 232 10039 2532 10139
rect 232 9883 2532 9983
rect 232 9727 2532 9827
rect 232 9571 2532 9671
rect 232 9415 2532 9515
rect 232 9259 2532 9359
rect 232 9103 2532 9203
rect 232 8947 2532 9047
rect 232 8791 2532 8891
rect 232 8635 2532 8735
rect 232 8479 2532 8579
rect 232 8323 2532 8423
rect 232 8167 2532 8267
rect 232 8011 2532 8111
rect 232 7855 2532 7955
rect 232 7699 2532 7799
rect 232 7543 2532 7643
rect 232 7387 2532 7487
rect 232 7231 2532 7331
rect 232 7075 2532 7175
rect 232 6919 2532 7019
rect 232 6763 2532 6863
rect 232 6607 2532 6707
rect 232 6451 2532 6551
rect 232 6295 2532 6395
rect 232 6139 2532 6239
rect 232 5983 2532 6083
rect 232 5827 2532 5927
rect 232 5671 2532 5771
rect 232 5515 2532 5615
rect 232 5359 2532 5459
rect 232 5203 2532 5303
rect 232 5047 2532 5147
rect 232 4891 2532 4991
rect 232 4735 2532 4835
rect 232 4579 2532 4679
rect 232 4423 2532 4523
rect 232 4267 2532 4367
rect 232 4111 2532 4211
rect 232 3955 2532 4055
rect 232 3799 2532 3899
rect 232 3643 2532 3743
rect 232 3487 2532 3587
rect 232 3331 2532 3431
rect 232 3175 2532 3275
rect 232 3019 2532 3119
rect 232 2863 2532 2963
rect 232 2707 2532 2807
rect 232 2551 2532 2651
rect 232 2395 2532 2495
rect 232 2239 2532 2339
rect 232 2083 2532 2183
rect 232 1927 2532 2027
rect 232 1771 2532 1871
rect 232 1615 2532 1715
rect 232 1459 2532 1559
rect 232 1303 2532 1403
rect 232 1147 2532 1247
rect 232 991 2532 1091
rect 232 835 2532 935
rect 232 679 2532 779
rect 232 523 2532 623
rect 232 367 2532 467
rect 232 211 2532 311
<< mvpdiff >>
rect 232 42944 2532 42956
rect 232 42910 240 42944
rect 2524 42910 2532 42944
rect 232 42899 2532 42910
rect 232 42788 2532 42799
rect 232 42754 240 42788
rect 2524 42754 2532 42788
rect 232 42743 2532 42754
rect 232 42632 2532 42643
rect 232 42598 240 42632
rect 2524 42598 2532 42632
rect 232 42587 2532 42598
rect 232 42476 2532 42487
rect 232 42442 240 42476
rect 2524 42442 2532 42476
rect 232 42431 2532 42442
rect 232 42320 2532 42331
rect 232 42286 240 42320
rect 2524 42286 2532 42320
rect 232 42275 2532 42286
rect 232 42164 2532 42175
rect 232 42130 240 42164
rect 2524 42130 2532 42164
rect 232 42119 2532 42130
rect 232 42008 2532 42019
rect 232 41974 240 42008
rect 2524 41974 2532 42008
rect 232 41963 2532 41974
rect 232 41852 2532 41863
rect 232 41818 240 41852
rect 2524 41818 2532 41852
rect 232 41807 2532 41818
rect 232 41696 2532 41707
rect 232 41662 240 41696
rect 2524 41662 2532 41696
rect 232 41651 2532 41662
rect 232 41540 2532 41551
rect 232 41506 240 41540
rect 2524 41506 2532 41540
rect 232 41495 2532 41506
rect 232 41384 2532 41395
rect 232 41350 240 41384
rect 2524 41350 2532 41384
rect 232 41339 2532 41350
rect 232 41228 2532 41239
rect 232 41194 240 41228
rect 2524 41194 2532 41228
rect 232 41183 2532 41194
rect 232 41072 2532 41083
rect 232 41038 240 41072
rect 2524 41038 2532 41072
rect 232 41027 2532 41038
rect 232 40916 2532 40927
rect 232 40882 240 40916
rect 2524 40882 2532 40916
rect 232 40871 2532 40882
rect 232 40760 2532 40771
rect 232 40726 240 40760
rect 2524 40726 2532 40760
rect 232 40715 2532 40726
rect 232 40604 2532 40615
rect 232 40570 240 40604
rect 2524 40570 2532 40604
rect 232 40559 2532 40570
rect 232 40448 2532 40459
rect 232 40414 240 40448
rect 2524 40414 2532 40448
rect 232 40403 2532 40414
rect 232 40292 2532 40303
rect 232 40258 240 40292
rect 2524 40258 2532 40292
rect 232 40247 2532 40258
rect 232 40136 2532 40147
rect 232 40102 240 40136
rect 2524 40102 2532 40136
rect 232 40091 2532 40102
rect 232 39980 2532 39991
rect 232 39946 240 39980
rect 2524 39946 2532 39980
rect 232 39935 2532 39946
rect 232 39824 2532 39835
rect 232 39790 240 39824
rect 2524 39790 2532 39824
rect 232 39779 2532 39790
rect 232 39668 2532 39679
rect 232 39634 240 39668
rect 2524 39634 2532 39668
rect 232 39623 2532 39634
rect 232 39512 2532 39523
rect 232 39478 240 39512
rect 2524 39478 2532 39512
rect 232 39467 2532 39478
rect 232 39356 2532 39367
rect 232 39322 240 39356
rect 2524 39322 2532 39356
rect 232 39311 2532 39322
rect 232 39200 2532 39211
rect 232 39166 240 39200
rect 2524 39166 2532 39200
rect 232 39155 2532 39166
rect 232 39044 2532 39055
rect 232 39010 240 39044
rect 2524 39010 2532 39044
rect 232 38999 2532 39010
rect 232 38888 2532 38899
rect 232 38854 240 38888
rect 2524 38854 2532 38888
rect 232 38843 2532 38854
rect 232 38732 2532 38743
rect 232 38698 240 38732
rect 2524 38698 2532 38732
rect 232 38687 2532 38698
rect 232 38576 2532 38587
rect 232 38542 240 38576
rect 2524 38542 2532 38576
rect 232 38531 2532 38542
rect 232 38420 2532 38431
rect 232 38386 240 38420
rect 2524 38386 2532 38420
rect 232 38375 2532 38386
rect 232 38264 2532 38275
rect 232 38230 240 38264
rect 2524 38230 2532 38264
rect 232 38219 2532 38230
rect 232 38108 2532 38119
rect 232 38074 240 38108
rect 2524 38074 2532 38108
rect 232 38063 2532 38074
rect 232 37952 2532 37963
rect 232 37918 240 37952
rect 2524 37918 2532 37952
rect 232 37907 2532 37918
rect 232 37796 2532 37807
rect 232 37762 240 37796
rect 2524 37762 2532 37796
rect 232 37751 2532 37762
rect 232 37640 2532 37651
rect 232 37606 240 37640
rect 2524 37606 2532 37640
rect 232 37595 2532 37606
rect 232 37484 2532 37495
rect 232 37450 240 37484
rect 2524 37450 2532 37484
rect 232 37439 2532 37450
rect 232 37328 2532 37339
rect 232 37294 240 37328
rect 2524 37294 2532 37328
rect 232 37283 2532 37294
rect 232 37172 2532 37183
rect 232 37138 240 37172
rect 2524 37138 2532 37172
rect 232 37127 2532 37138
rect 232 37016 2532 37027
rect 232 36982 240 37016
rect 2524 36982 2532 37016
rect 232 36971 2532 36982
rect 232 36860 2532 36871
rect 232 36826 240 36860
rect 2524 36826 2532 36860
rect 232 36815 2532 36826
rect 232 36704 2532 36715
rect 232 36670 240 36704
rect 2524 36670 2532 36704
rect 232 36659 2532 36670
rect 232 36548 2532 36559
rect 232 36514 240 36548
rect 2524 36514 2532 36548
rect 232 36503 2532 36514
rect 232 36392 2532 36403
rect 232 36358 240 36392
rect 2524 36358 2532 36392
rect 232 36347 2532 36358
rect 232 36236 2532 36247
rect 232 36202 240 36236
rect 2524 36202 2532 36236
rect 232 36191 2532 36202
rect 232 36080 2532 36091
rect 232 36046 240 36080
rect 2524 36046 2532 36080
rect 232 36035 2532 36046
rect 232 35924 2532 35935
rect 232 35890 240 35924
rect 2524 35890 2532 35924
rect 232 35879 2532 35890
rect 232 35768 2532 35779
rect 232 35734 240 35768
rect 2524 35734 2532 35768
rect 232 35723 2532 35734
rect 232 35612 2532 35623
rect 232 35578 240 35612
rect 2524 35578 2532 35612
rect 232 35567 2532 35578
rect 232 35456 2532 35467
rect 232 35422 240 35456
rect 2524 35422 2532 35456
rect 232 35411 2532 35422
rect 232 35300 2532 35311
rect 232 35266 240 35300
rect 2524 35266 2532 35300
rect 232 35255 2532 35266
rect 232 35144 2532 35155
rect 232 35110 240 35144
rect 2524 35110 2532 35144
rect 232 35099 2532 35110
rect 232 34988 2532 34999
rect 232 34954 240 34988
rect 2524 34954 2532 34988
rect 232 34943 2532 34954
rect 232 34832 2532 34843
rect 232 34798 240 34832
rect 2524 34798 2532 34832
rect 232 34787 2532 34798
rect 232 34676 2532 34687
rect 232 34642 240 34676
rect 2524 34642 2532 34676
rect 232 34631 2532 34642
rect 232 34520 2532 34531
rect 232 34486 240 34520
rect 2524 34486 2532 34520
rect 232 34475 2532 34486
rect 232 34364 2532 34375
rect 232 34330 240 34364
rect 2524 34330 2532 34364
rect 232 34319 2532 34330
rect 232 34208 2532 34219
rect 232 34174 240 34208
rect 2524 34174 2532 34208
rect 232 34163 2532 34174
rect 232 34052 2532 34063
rect 232 34018 240 34052
rect 2524 34018 2532 34052
rect 232 34007 2532 34018
rect 232 33896 2532 33907
rect 232 33862 240 33896
rect 2524 33862 2532 33896
rect 232 33851 2532 33862
rect 232 33740 2532 33751
rect 232 33706 240 33740
rect 2524 33706 2532 33740
rect 232 33695 2532 33706
rect 232 33584 2532 33595
rect 232 33550 240 33584
rect 2524 33550 2532 33584
rect 232 33539 2532 33550
rect 232 33428 2532 33439
rect 232 33394 240 33428
rect 2524 33394 2532 33428
rect 232 33383 2532 33394
rect 232 33272 2532 33283
rect 232 33238 240 33272
rect 2524 33238 2532 33272
rect 232 33227 2532 33238
rect 232 33116 2532 33127
rect 232 33082 240 33116
rect 2524 33082 2532 33116
rect 232 33071 2532 33082
rect 232 32960 2532 32971
rect 232 32926 240 32960
rect 2524 32926 2532 32960
rect 232 32915 2532 32926
rect 232 32804 2532 32815
rect 232 32770 240 32804
rect 2524 32770 2532 32804
rect 232 32759 2532 32770
rect 232 32648 2532 32659
rect 232 32614 240 32648
rect 2524 32614 2532 32648
rect 232 32603 2532 32614
rect 232 32492 2532 32503
rect 232 32458 240 32492
rect 2524 32458 2532 32492
rect 232 32447 2532 32458
rect 232 32336 2532 32347
rect 232 32302 240 32336
rect 2524 32302 2532 32336
rect 232 32291 2532 32302
rect 232 32180 2532 32191
rect 232 32146 240 32180
rect 2524 32146 2532 32180
rect 232 32135 2532 32146
rect 232 32024 2532 32035
rect 232 31990 240 32024
rect 2524 31990 2532 32024
rect 232 31979 2532 31990
rect 232 31868 2532 31879
rect 232 31834 240 31868
rect 2524 31834 2532 31868
rect 232 31823 2532 31834
rect 232 31712 2532 31723
rect 232 31678 240 31712
rect 2524 31678 2532 31712
rect 232 31667 2532 31678
rect 232 31556 2532 31567
rect 232 31522 240 31556
rect 2524 31522 2532 31556
rect 232 31511 2532 31522
rect 232 31400 2532 31411
rect 232 31366 240 31400
rect 2524 31366 2532 31400
rect 232 31355 2532 31366
rect 232 31244 2532 31255
rect 232 31210 240 31244
rect 2524 31210 2532 31244
rect 232 31199 2532 31210
rect 232 31088 2532 31099
rect 232 31054 240 31088
rect 2524 31054 2532 31088
rect 232 31043 2532 31054
rect 232 30932 2532 30943
rect 232 30898 240 30932
rect 2524 30898 2532 30932
rect 232 30887 2532 30898
rect 232 30776 2532 30787
rect 232 30742 240 30776
rect 2524 30742 2532 30776
rect 232 30731 2532 30742
rect 232 30620 2532 30631
rect 232 30586 240 30620
rect 2524 30586 2532 30620
rect 232 30575 2532 30586
rect 232 30464 2532 30475
rect 232 30430 240 30464
rect 2524 30430 2532 30464
rect 232 30419 2532 30430
rect 232 30308 2532 30319
rect 232 30274 240 30308
rect 2524 30274 2532 30308
rect 232 30263 2532 30274
rect 232 30152 2532 30163
rect 232 30118 240 30152
rect 2524 30118 2532 30152
rect 232 30107 2532 30118
rect 232 29996 2532 30007
rect 232 29962 240 29996
rect 2524 29962 2532 29996
rect 232 29951 2532 29962
rect 232 29840 2532 29851
rect 232 29806 240 29840
rect 2524 29806 2532 29840
rect 232 29795 2532 29806
rect 232 29684 2532 29695
rect 232 29650 240 29684
rect 2524 29650 2532 29684
rect 232 29639 2532 29650
rect 232 29528 2532 29539
rect 232 29494 240 29528
rect 2524 29494 2532 29528
rect 232 29483 2532 29494
rect 232 29372 2532 29383
rect 232 29338 240 29372
rect 2524 29338 2532 29372
rect 232 29327 2532 29338
rect 232 29216 2532 29227
rect 232 29182 240 29216
rect 2524 29182 2532 29216
rect 232 29171 2532 29182
rect 232 29060 2532 29071
rect 232 29026 240 29060
rect 2524 29026 2532 29060
rect 232 29015 2532 29026
rect 232 28904 2532 28915
rect 232 28870 240 28904
rect 2524 28870 2532 28904
rect 232 28859 2532 28870
rect 232 28748 2532 28759
rect 232 28714 240 28748
rect 2524 28714 2532 28748
rect 232 28703 2532 28714
rect 232 28592 2532 28603
rect 232 28558 240 28592
rect 2524 28558 2532 28592
rect 232 28547 2532 28558
rect 232 28436 2532 28447
rect 232 28402 240 28436
rect 2524 28402 2532 28436
rect 232 28391 2532 28402
rect 232 28280 2532 28291
rect 232 28246 240 28280
rect 2524 28246 2532 28280
rect 232 28235 2532 28246
rect 232 28124 2532 28135
rect 232 28090 240 28124
rect 2524 28090 2532 28124
rect 232 28079 2532 28090
rect 232 27968 2532 27979
rect 232 27934 240 27968
rect 2524 27934 2532 27968
rect 232 27923 2532 27934
rect 232 27812 2532 27823
rect 232 27778 240 27812
rect 2524 27778 2532 27812
rect 232 27767 2532 27778
rect 232 27656 2532 27667
rect 232 27622 240 27656
rect 2524 27622 2532 27656
rect 232 27611 2532 27622
rect 232 27500 2532 27511
rect 232 27466 240 27500
rect 2524 27466 2532 27500
rect 232 27455 2532 27466
rect 232 27344 2532 27355
rect 232 27310 240 27344
rect 2524 27310 2532 27344
rect 232 27299 2532 27310
rect 232 27188 2532 27199
rect 232 27154 240 27188
rect 2524 27154 2532 27188
rect 232 27143 2532 27154
rect 232 27032 2532 27043
rect 232 26998 240 27032
rect 2524 26998 2532 27032
rect 232 26987 2532 26998
rect 232 26876 2532 26887
rect 232 26842 240 26876
rect 2524 26842 2532 26876
rect 232 26831 2532 26842
rect 232 26720 2532 26731
rect 232 26686 240 26720
rect 2524 26686 2532 26720
rect 232 26675 2532 26686
rect 232 26564 2532 26575
rect 232 26530 240 26564
rect 2524 26530 2532 26564
rect 232 26519 2532 26530
rect 232 26408 2532 26419
rect 232 26374 240 26408
rect 2524 26374 2532 26408
rect 232 26363 2532 26374
rect 232 26252 2532 26263
rect 232 26218 240 26252
rect 2524 26218 2532 26252
rect 232 26207 2532 26218
rect 232 26096 2532 26107
rect 232 26062 240 26096
rect 2524 26062 2532 26096
rect 232 26051 2532 26062
rect 232 25940 2532 25951
rect 232 25906 240 25940
rect 2524 25906 2532 25940
rect 232 25895 2532 25906
rect 232 25784 2532 25795
rect 232 25750 240 25784
rect 2524 25750 2532 25784
rect 232 25739 2532 25750
rect 232 25628 2532 25639
rect 232 25594 240 25628
rect 2524 25594 2532 25628
rect 232 25583 2532 25594
rect 232 25472 2532 25483
rect 232 25438 240 25472
rect 2524 25438 2532 25472
rect 232 25427 2532 25438
rect 232 25316 2532 25327
rect 232 25282 240 25316
rect 2524 25282 2532 25316
rect 232 25271 2532 25282
rect 232 25160 2532 25171
rect 232 25126 240 25160
rect 2524 25126 2532 25160
rect 232 25115 2532 25126
rect 232 25004 2532 25015
rect 232 24970 240 25004
rect 2524 24970 2532 25004
rect 232 24959 2532 24970
rect 232 24848 2532 24859
rect 232 24814 240 24848
rect 2524 24814 2532 24848
rect 232 24803 2532 24814
rect 232 24692 2532 24703
rect 232 24658 240 24692
rect 2524 24658 2532 24692
rect 232 24647 2532 24658
rect 232 24536 2532 24547
rect 232 24502 240 24536
rect 2524 24502 2532 24536
rect 232 24491 2532 24502
rect 232 24380 2532 24391
rect 232 24346 240 24380
rect 2524 24346 2532 24380
rect 232 24335 2532 24346
rect 232 24224 2532 24235
rect 232 24190 240 24224
rect 2524 24190 2532 24224
rect 232 24179 2532 24190
rect 232 24068 2532 24079
rect 232 24034 240 24068
rect 2524 24034 2532 24068
rect 232 24023 2532 24034
rect 232 23912 2532 23923
rect 232 23878 240 23912
rect 2524 23878 2532 23912
rect 232 23867 2532 23878
rect 232 23756 2532 23767
rect 232 23722 240 23756
rect 2524 23722 2532 23756
rect 232 23711 2532 23722
rect 232 23600 2532 23611
rect 232 23566 240 23600
rect 2524 23566 2532 23600
rect 232 23555 2532 23566
rect 232 23444 2532 23455
rect 232 23410 240 23444
rect 2524 23410 2532 23444
rect 232 23399 2532 23410
rect 232 23288 2532 23299
rect 232 23254 240 23288
rect 2524 23254 2532 23288
rect 232 23243 2532 23254
rect 232 23132 2532 23143
rect 232 23098 240 23132
rect 2524 23098 2532 23132
rect 232 23087 2532 23098
rect 232 22976 2532 22987
rect 232 22942 240 22976
rect 2524 22942 2532 22976
rect 232 22931 2532 22942
rect 232 22820 2532 22831
rect 232 22786 240 22820
rect 2524 22786 2532 22820
rect 232 22775 2532 22786
rect 232 22664 2532 22675
rect 232 22630 240 22664
rect 2524 22630 2532 22664
rect 232 22619 2532 22630
rect 232 22508 2532 22519
rect 232 22474 240 22508
rect 2524 22474 2532 22508
rect 232 22463 2532 22474
rect 232 22352 2532 22363
rect 232 22318 240 22352
rect 2524 22318 2532 22352
rect 232 22307 2532 22318
rect 232 22196 2532 22207
rect 232 22162 240 22196
rect 2524 22162 2532 22196
rect 232 22151 2532 22162
rect 232 22040 2532 22051
rect 232 22006 240 22040
rect 2524 22006 2532 22040
rect 232 21995 2532 22006
rect 232 21884 2532 21895
rect 232 21850 240 21884
rect 2524 21850 2532 21884
rect 232 21839 2532 21850
rect 232 21728 2532 21739
rect 232 21694 240 21728
rect 2524 21694 2532 21728
rect 232 21683 2532 21694
rect 232 21572 2532 21583
rect 232 21538 240 21572
rect 2524 21538 2532 21572
rect 232 21527 2532 21538
rect 232 21416 2532 21427
rect 232 21382 240 21416
rect 2524 21382 2532 21416
rect 232 21371 2532 21382
rect 232 21260 2532 21271
rect 232 21226 240 21260
rect 2524 21226 2532 21260
rect 232 21215 2532 21226
rect 232 21104 2532 21115
rect 232 21070 240 21104
rect 2524 21070 2532 21104
rect 232 21059 2532 21070
rect 232 20948 2532 20959
rect 232 20914 240 20948
rect 2524 20914 2532 20948
rect 232 20903 2532 20914
rect 232 20792 2532 20803
rect 232 20758 240 20792
rect 2524 20758 2532 20792
rect 232 20747 2532 20758
rect 232 20636 2532 20647
rect 232 20602 240 20636
rect 2524 20602 2532 20636
rect 232 20591 2532 20602
rect 232 20480 2532 20491
rect 232 20446 240 20480
rect 2524 20446 2532 20480
rect 232 20435 2532 20446
rect 232 20324 2532 20335
rect 232 20290 240 20324
rect 2524 20290 2532 20324
rect 232 20279 2532 20290
rect 232 20168 2532 20179
rect 232 20134 240 20168
rect 2524 20134 2532 20168
rect 232 20123 2532 20134
rect 232 20012 2532 20023
rect 232 19978 240 20012
rect 2524 19978 2532 20012
rect 232 19967 2532 19978
rect 232 19856 2532 19867
rect 232 19822 240 19856
rect 2524 19822 2532 19856
rect 232 19811 2532 19822
rect 232 19700 2532 19711
rect 232 19666 240 19700
rect 2524 19666 2532 19700
rect 232 19655 2532 19666
rect 232 19544 2532 19555
rect 232 19510 240 19544
rect 2524 19510 2532 19544
rect 232 19499 2532 19510
rect 232 19388 2532 19399
rect 232 19354 240 19388
rect 2524 19354 2532 19388
rect 232 19343 2532 19354
rect 232 19232 2532 19243
rect 232 19198 240 19232
rect 2524 19198 2532 19232
rect 232 19187 2532 19198
rect 232 19076 2532 19087
rect 232 19042 240 19076
rect 2524 19042 2532 19076
rect 232 19031 2532 19042
rect 232 18920 2532 18931
rect 232 18886 240 18920
rect 2524 18886 2532 18920
rect 232 18875 2532 18886
rect 232 18764 2532 18775
rect 232 18730 240 18764
rect 2524 18730 2532 18764
rect 232 18719 2532 18730
rect 232 18608 2532 18619
rect 232 18574 240 18608
rect 2524 18574 2532 18608
rect 232 18563 2532 18574
rect 232 18452 2532 18463
rect 232 18418 240 18452
rect 2524 18418 2532 18452
rect 232 18407 2532 18418
rect 232 18296 2532 18307
rect 232 18262 240 18296
rect 2524 18262 2532 18296
rect 232 18251 2532 18262
rect 232 18140 2532 18151
rect 232 18106 240 18140
rect 2524 18106 2532 18140
rect 232 18095 2532 18106
rect 232 17984 2532 17995
rect 232 17950 240 17984
rect 2524 17950 2532 17984
rect 232 17939 2532 17950
rect 232 17828 2532 17839
rect 232 17794 240 17828
rect 2524 17794 2532 17828
rect 232 17783 2532 17794
rect 232 17672 2532 17683
rect 232 17638 240 17672
rect 2524 17638 2532 17672
rect 232 17627 2532 17638
rect 232 17516 2532 17527
rect 232 17482 240 17516
rect 2524 17482 2532 17516
rect 232 17471 2532 17482
rect 232 17360 2532 17371
rect 232 17326 240 17360
rect 2524 17326 2532 17360
rect 232 17315 2532 17326
rect 232 17204 2532 17215
rect 232 17170 240 17204
rect 2524 17170 2532 17204
rect 232 17159 2532 17170
rect 232 17048 2532 17059
rect 232 17014 240 17048
rect 2524 17014 2532 17048
rect 232 17003 2532 17014
rect 232 16892 2532 16903
rect 232 16858 240 16892
rect 2524 16858 2532 16892
rect 232 16847 2532 16858
rect 232 16736 2532 16747
rect 232 16702 240 16736
rect 2524 16702 2532 16736
rect 232 16691 2532 16702
rect 232 16580 2532 16591
rect 232 16546 240 16580
rect 2524 16546 2532 16580
rect 232 16535 2532 16546
rect 232 16424 2532 16435
rect 232 16390 240 16424
rect 2524 16390 2532 16424
rect 232 16379 2532 16390
rect 232 16268 2532 16279
rect 232 16234 240 16268
rect 2524 16234 2532 16268
rect 232 16223 2532 16234
rect 232 16112 2532 16123
rect 232 16078 240 16112
rect 2524 16078 2532 16112
rect 232 16067 2532 16078
rect 232 15956 2532 15967
rect 232 15922 240 15956
rect 2524 15922 2532 15956
rect 232 15911 2532 15922
rect 232 15800 2532 15811
rect 232 15766 240 15800
rect 2524 15766 2532 15800
rect 232 15755 2532 15766
rect 232 15644 2532 15655
rect 232 15610 240 15644
rect 2524 15610 2532 15644
rect 232 15599 2532 15610
rect 232 15488 2532 15499
rect 232 15454 240 15488
rect 2524 15454 2532 15488
rect 232 15443 2532 15454
rect 232 15332 2532 15343
rect 232 15298 240 15332
rect 2524 15298 2532 15332
rect 232 15287 2532 15298
rect 232 15176 2532 15187
rect 232 15142 240 15176
rect 2524 15142 2532 15176
rect 232 15131 2532 15142
rect 232 15020 2532 15031
rect 232 14986 240 15020
rect 2524 14986 2532 15020
rect 232 14975 2532 14986
rect 232 14864 2532 14875
rect 232 14830 240 14864
rect 2524 14830 2532 14864
rect 232 14819 2532 14830
rect 232 14708 2532 14719
rect 232 14674 240 14708
rect 2524 14674 2532 14708
rect 232 14663 2532 14674
rect 232 14552 2532 14563
rect 232 14518 240 14552
rect 2524 14518 2532 14552
rect 232 14507 2532 14518
rect 232 14396 2532 14407
rect 232 14362 240 14396
rect 2524 14362 2532 14396
rect 232 14351 2532 14362
rect 232 14240 2532 14251
rect 232 14206 240 14240
rect 2524 14206 2532 14240
rect 232 14195 2532 14206
rect 232 14084 2532 14095
rect 232 14050 240 14084
rect 2524 14050 2532 14084
rect 232 14039 2532 14050
rect 232 13928 2532 13939
rect 232 13894 240 13928
rect 2524 13894 2532 13928
rect 232 13883 2532 13894
rect 232 13772 2532 13783
rect 232 13738 240 13772
rect 2524 13738 2532 13772
rect 232 13727 2532 13738
rect 232 13616 2532 13627
rect 232 13582 240 13616
rect 2524 13582 2532 13616
rect 232 13571 2532 13582
rect 232 13460 2532 13471
rect 232 13426 240 13460
rect 2524 13426 2532 13460
rect 232 13415 2532 13426
rect 232 13304 2532 13315
rect 232 13270 240 13304
rect 2524 13270 2532 13304
rect 232 13259 2532 13270
rect 232 13148 2532 13159
rect 232 13114 240 13148
rect 2524 13114 2532 13148
rect 232 13103 2532 13114
rect 232 12992 2532 13003
rect 232 12958 240 12992
rect 2524 12958 2532 12992
rect 232 12947 2532 12958
rect 232 12836 2532 12847
rect 232 12802 240 12836
rect 2524 12802 2532 12836
rect 232 12791 2532 12802
rect 232 12680 2532 12691
rect 232 12646 240 12680
rect 2524 12646 2532 12680
rect 232 12635 2532 12646
rect 232 12524 2532 12535
rect 232 12490 240 12524
rect 2524 12490 2532 12524
rect 232 12479 2532 12490
rect 232 12368 2532 12379
rect 232 12334 240 12368
rect 2524 12334 2532 12368
rect 232 12323 2532 12334
rect 232 12212 2532 12223
rect 232 12178 240 12212
rect 2524 12178 2532 12212
rect 232 12167 2532 12178
rect 232 12056 2532 12067
rect 232 12022 240 12056
rect 2524 12022 2532 12056
rect 232 12011 2532 12022
rect 232 11900 2532 11911
rect 232 11866 240 11900
rect 2524 11866 2532 11900
rect 232 11855 2532 11866
rect 232 11744 2532 11755
rect 232 11710 240 11744
rect 2524 11710 2532 11744
rect 232 11699 2532 11710
rect 232 11588 2532 11599
rect 232 11554 240 11588
rect 2524 11554 2532 11588
rect 232 11543 2532 11554
rect 232 11432 2532 11443
rect 232 11398 240 11432
rect 2524 11398 2532 11432
rect 232 11387 2532 11398
rect 232 11276 2532 11287
rect 232 11242 240 11276
rect 2524 11242 2532 11276
rect 232 11231 2532 11242
rect 232 11120 2532 11131
rect 232 11086 240 11120
rect 2524 11086 2532 11120
rect 232 11075 2532 11086
rect 232 10964 2532 10975
rect 232 10930 240 10964
rect 2524 10930 2532 10964
rect 232 10919 2532 10930
rect 232 10808 2532 10819
rect 232 10774 240 10808
rect 2524 10774 2532 10808
rect 232 10763 2532 10774
rect 232 10652 2532 10663
rect 232 10618 240 10652
rect 2524 10618 2532 10652
rect 232 10607 2532 10618
rect 232 10496 2532 10507
rect 232 10462 240 10496
rect 2524 10462 2532 10496
rect 232 10451 2532 10462
rect 232 10340 2532 10351
rect 232 10306 240 10340
rect 2524 10306 2532 10340
rect 232 10295 2532 10306
rect 232 10184 2532 10195
rect 232 10150 240 10184
rect 2524 10150 2532 10184
rect 232 10139 2532 10150
rect 232 10028 2532 10039
rect 232 9994 240 10028
rect 2524 9994 2532 10028
rect 232 9983 2532 9994
rect 232 9872 2532 9883
rect 232 9838 240 9872
rect 2524 9838 2532 9872
rect 232 9827 2532 9838
rect 232 9716 2532 9727
rect 232 9682 240 9716
rect 2524 9682 2532 9716
rect 232 9671 2532 9682
rect 232 9560 2532 9571
rect 232 9526 240 9560
rect 2524 9526 2532 9560
rect 232 9515 2532 9526
rect 232 9404 2532 9415
rect 232 9370 240 9404
rect 2524 9370 2532 9404
rect 232 9359 2532 9370
rect 232 9248 2532 9259
rect 232 9214 240 9248
rect 2524 9214 2532 9248
rect 232 9203 2532 9214
rect 232 9092 2532 9103
rect 232 9058 240 9092
rect 2524 9058 2532 9092
rect 232 9047 2532 9058
rect 232 8936 2532 8947
rect 232 8902 240 8936
rect 2524 8902 2532 8936
rect 232 8891 2532 8902
rect 232 8780 2532 8791
rect 232 8746 240 8780
rect 2524 8746 2532 8780
rect 232 8735 2532 8746
rect 232 8624 2532 8635
rect 232 8590 240 8624
rect 2524 8590 2532 8624
rect 232 8579 2532 8590
rect 232 8468 2532 8479
rect 232 8434 240 8468
rect 2524 8434 2532 8468
rect 232 8423 2532 8434
rect 232 8312 2532 8323
rect 232 8278 240 8312
rect 2524 8278 2532 8312
rect 232 8267 2532 8278
rect 232 8156 2532 8167
rect 232 8122 240 8156
rect 2524 8122 2532 8156
rect 232 8111 2532 8122
rect 232 8000 2532 8011
rect 232 7966 240 8000
rect 2524 7966 2532 8000
rect 232 7955 2532 7966
rect 232 7844 2532 7855
rect 232 7810 240 7844
rect 2524 7810 2532 7844
rect 232 7799 2532 7810
rect 232 7688 2532 7699
rect 232 7654 240 7688
rect 2524 7654 2532 7688
rect 232 7643 2532 7654
rect 232 7532 2532 7543
rect 232 7498 240 7532
rect 2524 7498 2532 7532
rect 232 7487 2532 7498
rect 232 7376 2532 7387
rect 232 7342 240 7376
rect 2524 7342 2532 7376
rect 232 7331 2532 7342
rect 232 7220 2532 7231
rect 232 7186 240 7220
rect 2524 7186 2532 7220
rect 232 7175 2532 7186
rect 232 7064 2532 7075
rect 232 7030 240 7064
rect 2524 7030 2532 7064
rect 232 7019 2532 7030
rect 232 6908 2532 6919
rect 232 6874 240 6908
rect 2524 6874 2532 6908
rect 232 6863 2532 6874
rect 232 6752 2532 6763
rect 232 6718 240 6752
rect 2524 6718 2532 6752
rect 232 6707 2532 6718
rect 232 6596 2532 6607
rect 232 6562 240 6596
rect 2524 6562 2532 6596
rect 232 6551 2532 6562
rect 232 6440 2532 6451
rect 232 6406 240 6440
rect 2524 6406 2532 6440
rect 232 6395 2532 6406
rect 232 6284 2532 6295
rect 232 6250 240 6284
rect 2524 6250 2532 6284
rect 232 6239 2532 6250
rect 232 6128 2532 6139
rect 232 6094 240 6128
rect 2524 6094 2532 6128
rect 232 6083 2532 6094
rect 232 5972 2532 5983
rect 232 5938 240 5972
rect 2524 5938 2532 5972
rect 232 5927 2532 5938
rect 232 5816 2532 5827
rect 232 5782 240 5816
rect 2524 5782 2532 5816
rect 232 5771 2532 5782
rect 232 5660 2532 5671
rect 232 5626 240 5660
rect 2524 5626 2532 5660
rect 232 5615 2532 5626
rect 232 5504 2532 5515
rect 232 5470 240 5504
rect 2524 5470 2532 5504
rect 232 5459 2532 5470
rect 232 5348 2532 5359
rect 232 5314 240 5348
rect 2524 5314 2532 5348
rect 232 5303 2532 5314
rect 232 5192 2532 5203
rect 232 5158 240 5192
rect 2524 5158 2532 5192
rect 232 5147 2532 5158
rect 232 5036 2532 5047
rect 232 5002 240 5036
rect 2524 5002 2532 5036
rect 232 4991 2532 5002
rect 232 4880 2532 4891
rect 232 4846 240 4880
rect 2524 4846 2532 4880
rect 232 4835 2532 4846
rect 232 4724 2532 4735
rect 232 4690 240 4724
rect 2524 4690 2532 4724
rect 232 4679 2532 4690
rect 232 4568 2532 4579
rect 232 4534 240 4568
rect 2524 4534 2532 4568
rect 232 4523 2532 4534
rect 232 4412 2532 4423
rect 232 4378 240 4412
rect 2524 4378 2532 4412
rect 232 4367 2532 4378
rect 232 4256 2532 4267
rect 232 4222 240 4256
rect 2524 4222 2532 4256
rect 232 4211 2532 4222
rect 232 4100 2532 4111
rect 232 4066 240 4100
rect 2524 4066 2532 4100
rect 232 4055 2532 4066
rect 232 3944 2532 3955
rect 232 3910 240 3944
rect 2524 3910 2532 3944
rect 232 3899 2532 3910
rect 232 3788 2532 3799
rect 232 3754 240 3788
rect 2524 3754 2532 3788
rect 232 3743 2532 3754
rect 232 3632 2532 3643
rect 232 3598 240 3632
rect 2524 3598 2532 3632
rect 232 3587 2532 3598
rect 232 3476 2532 3487
rect 232 3442 240 3476
rect 2524 3442 2532 3476
rect 232 3431 2532 3442
rect 232 3320 2532 3331
rect 232 3286 240 3320
rect 2524 3286 2532 3320
rect 232 3275 2532 3286
rect 232 3164 2532 3175
rect 232 3130 240 3164
rect 2524 3130 2532 3164
rect 232 3119 2532 3130
rect 232 3008 2532 3019
rect 232 2974 240 3008
rect 2524 2974 2532 3008
rect 232 2963 2532 2974
rect 232 2852 2532 2863
rect 232 2818 240 2852
rect 2524 2818 2532 2852
rect 232 2807 2532 2818
rect 232 2696 2532 2707
rect 232 2662 240 2696
rect 2524 2662 2532 2696
rect 232 2651 2532 2662
rect 232 2540 2532 2551
rect 232 2506 240 2540
rect 2524 2506 2532 2540
rect 232 2495 2532 2506
rect 232 2384 2532 2395
rect 232 2350 240 2384
rect 2524 2350 2532 2384
rect 232 2339 2532 2350
rect 232 2228 2532 2239
rect 232 2194 240 2228
rect 2524 2194 2532 2228
rect 232 2183 2532 2194
rect 232 2072 2532 2083
rect 232 2038 240 2072
rect 2524 2038 2532 2072
rect 232 2027 2532 2038
rect 232 1916 2532 1927
rect 232 1882 240 1916
rect 2524 1882 2532 1916
rect 232 1871 2532 1882
rect 232 1760 2532 1771
rect 232 1726 240 1760
rect 2524 1726 2532 1760
rect 232 1715 2532 1726
rect 232 1604 2532 1615
rect 232 1570 240 1604
rect 2524 1570 2532 1604
rect 232 1559 2532 1570
rect 232 1448 2532 1459
rect 232 1414 240 1448
rect 2524 1414 2532 1448
rect 232 1403 2532 1414
rect 232 1292 2532 1303
rect 232 1258 240 1292
rect 2524 1258 2532 1292
rect 232 1247 2532 1258
rect 232 1136 2532 1147
rect 232 1102 240 1136
rect 2524 1102 2532 1136
rect 232 1091 2532 1102
rect 232 980 2532 991
rect 232 946 240 980
rect 2524 946 2532 980
rect 232 935 2532 946
rect 232 824 2532 835
rect 232 790 240 824
rect 2524 790 2532 824
rect 232 779 2532 790
rect 232 668 2532 679
rect 232 634 240 668
rect 2524 634 2532 668
rect 232 623 2532 634
rect 232 512 2532 523
rect 232 478 240 512
rect 2524 478 2532 512
rect 232 467 2532 478
rect 232 356 2532 367
rect 232 322 240 356
rect 2524 322 2532 356
rect 232 311 2532 322
rect 232 200 2532 211
rect 232 166 240 200
rect 2524 166 2532 200
rect 232 154 2532 166
<< mvpdiffc >>
rect 240 42910 2524 42944
rect 240 42754 2524 42788
rect 240 42598 2524 42632
rect 240 42442 2524 42476
rect 240 42286 2524 42320
rect 240 42130 2524 42164
rect 240 41974 2524 42008
rect 240 41818 2524 41852
rect 240 41662 2524 41696
rect 240 41506 2524 41540
rect 240 41350 2524 41384
rect 240 41194 2524 41228
rect 240 41038 2524 41072
rect 240 40882 2524 40916
rect 240 40726 2524 40760
rect 240 40570 2524 40604
rect 240 40414 2524 40448
rect 240 40258 2524 40292
rect 240 40102 2524 40136
rect 240 39946 2524 39980
rect 240 39790 2524 39824
rect 240 39634 2524 39668
rect 240 39478 2524 39512
rect 240 39322 2524 39356
rect 240 39166 2524 39200
rect 240 39010 2524 39044
rect 240 38854 2524 38888
rect 240 38698 2524 38732
rect 240 38542 2524 38576
rect 240 38386 2524 38420
rect 240 38230 2524 38264
rect 240 38074 2524 38108
rect 240 37918 2524 37952
rect 240 37762 2524 37796
rect 240 37606 2524 37640
rect 240 37450 2524 37484
rect 240 37294 2524 37328
rect 240 37138 2524 37172
rect 240 36982 2524 37016
rect 240 36826 2524 36860
rect 240 36670 2524 36704
rect 240 36514 2524 36548
rect 240 36358 2524 36392
rect 240 36202 2524 36236
rect 240 36046 2524 36080
rect 240 35890 2524 35924
rect 240 35734 2524 35768
rect 240 35578 2524 35612
rect 240 35422 2524 35456
rect 240 35266 2524 35300
rect 240 35110 2524 35144
rect 240 34954 2524 34988
rect 240 34798 2524 34832
rect 240 34642 2524 34676
rect 240 34486 2524 34520
rect 240 34330 2524 34364
rect 240 34174 2524 34208
rect 240 34018 2524 34052
rect 240 33862 2524 33896
rect 240 33706 2524 33740
rect 240 33550 2524 33584
rect 240 33394 2524 33428
rect 240 33238 2524 33272
rect 240 33082 2524 33116
rect 240 32926 2524 32960
rect 240 32770 2524 32804
rect 240 32614 2524 32648
rect 240 32458 2524 32492
rect 240 32302 2524 32336
rect 240 32146 2524 32180
rect 240 31990 2524 32024
rect 240 31834 2524 31868
rect 240 31678 2524 31712
rect 240 31522 2524 31556
rect 240 31366 2524 31400
rect 240 31210 2524 31244
rect 240 31054 2524 31088
rect 240 30898 2524 30932
rect 240 30742 2524 30776
rect 240 30586 2524 30620
rect 240 30430 2524 30464
rect 240 30274 2524 30308
rect 240 30118 2524 30152
rect 240 29962 2524 29996
rect 240 29806 2524 29840
rect 240 29650 2524 29684
rect 240 29494 2524 29528
rect 240 29338 2524 29372
rect 240 29182 2524 29216
rect 240 29026 2524 29060
rect 240 28870 2524 28904
rect 240 28714 2524 28748
rect 240 28558 2524 28592
rect 240 28402 2524 28436
rect 240 28246 2524 28280
rect 240 28090 2524 28124
rect 240 27934 2524 27968
rect 240 27778 2524 27812
rect 240 27622 2524 27656
rect 240 27466 2524 27500
rect 240 27310 2524 27344
rect 240 27154 2524 27188
rect 240 26998 2524 27032
rect 240 26842 2524 26876
rect 240 26686 2524 26720
rect 240 26530 2524 26564
rect 240 26374 2524 26408
rect 240 26218 2524 26252
rect 240 26062 2524 26096
rect 240 25906 2524 25940
rect 240 25750 2524 25784
rect 240 25594 2524 25628
rect 240 25438 2524 25472
rect 240 25282 2524 25316
rect 240 25126 2524 25160
rect 240 24970 2524 25004
rect 240 24814 2524 24848
rect 240 24658 2524 24692
rect 240 24502 2524 24536
rect 240 24346 2524 24380
rect 240 24190 2524 24224
rect 240 24034 2524 24068
rect 240 23878 2524 23912
rect 240 23722 2524 23756
rect 240 23566 2524 23600
rect 240 23410 2524 23444
rect 240 23254 2524 23288
rect 240 23098 2524 23132
rect 240 22942 2524 22976
rect 240 22786 2524 22820
rect 240 22630 2524 22664
rect 240 22474 2524 22508
rect 240 22318 2524 22352
rect 240 22162 2524 22196
rect 240 22006 2524 22040
rect 240 21850 2524 21884
rect 240 21694 2524 21728
rect 240 21538 2524 21572
rect 240 21382 2524 21416
rect 240 21226 2524 21260
rect 240 21070 2524 21104
rect 240 20914 2524 20948
rect 240 20758 2524 20792
rect 240 20602 2524 20636
rect 240 20446 2524 20480
rect 240 20290 2524 20324
rect 240 20134 2524 20168
rect 240 19978 2524 20012
rect 240 19822 2524 19856
rect 240 19666 2524 19700
rect 240 19510 2524 19544
rect 240 19354 2524 19388
rect 240 19198 2524 19232
rect 240 19042 2524 19076
rect 240 18886 2524 18920
rect 240 18730 2524 18764
rect 240 18574 2524 18608
rect 240 18418 2524 18452
rect 240 18262 2524 18296
rect 240 18106 2524 18140
rect 240 17950 2524 17984
rect 240 17794 2524 17828
rect 240 17638 2524 17672
rect 240 17482 2524 17516
rect 240 17326 2524 17360
rect 240 17170 2524 17204
rect 240 17014 2524 17048
rect 240 16858 2524 16892
rect 240 16702 2524 16736
rect 240 16546 2524 16580
rect 240 16390 2524 16424
rect 240 16234 2524 16268
rect 240 16078 2524 16112
rect 240 15922 2524 15956
rect 240 15766 2524 15800
rect 240 15610 2524 15644
rect 240 15454 2524 15488
rect 240 15298 2524 15332
rect 240 15142 2524 15176
rect 240 14986 2524 15020
rect 240 14830 2524 14864
rect 240 14674 2524 14708
rect 240 14518 2524 14552
rect 240 14362 2524 14396
rect 240 14206 2524 14240
rect 240 14050 2524 14084
rect 240 13894 2524 13928
rect 240 13738 2524 13772
rect 240 13582 2524 13616
rect 240 13426 2524 13460
rect 240 13270 2524 13304
rect 240 13114 2524 13148
rect 240 12958 2524 12992
rect 240 12802 2524 12836
rect 240 12646 2524 12680
rect 240 12490 2524 12524
rect 240 12334 2524 12368
rect 240 12178 2524 12212
rect 240 12022 2524 12056
rect 240 11866 2524 11900
rect 240 11710 2524 11744
rect 240 11554 2524 11588
rect 240 11398 2524 11432
rect 240 11242 2524 11276
rect 240 11086 2524 11120
rect 240 10930 2524 10964
rect 240 10774 2524 10808
rect 240 10618 2524 10652
rect 240 10462 2524 10496
rect 240 10306 2524 10340
rect 240 10150 2524 10184
rect 240 9994 2524 10028
rect 240 9838 2524 9872
rect 240 9682 2524 9716
rect 240 9526 2524 9560
rect 240 9370 2524 9404
rect 240 9214 2524 9248
rect 240 9058 2524 9092
rect 240 8902 2524 8936
rect 240 8746 2524 8780
rect 240 8590 2524 8624
rect 240 8434 2524 8468
rect 240 8278 2524 8312
rect 240 8122 2524 8156
rect 240 7966 2524 8000
rect 240 7810 2524 7844
rect 240 7654 2524 7688
rect 240 7498 2524 7532
rect 240 7342 2524 7376
rect 240 7186 2524 7220
rect 240 7030 2524 7064
rect 240 6874 2524 6908
rect 240 6718 2524 6752
rect 240 6562 2524 6596
rect 240 6406 2524 6440
rect 240 6250 2524 6284
rect 240 6094 2524 6128
rect 240 5938 2524 5972
rect 240 5782 2524 5816
rect 240 5626 2524 5660
rect 240 5470 2524 5504
rect 240 5314 2524 5348
rect 240 5158 2524 5192
rect 240 5002 2524 5036
rect 240 4846 2524 4880
rect 240 4690 2524 4724
rect 240 4534 2524 4568
rect 240 4378 2524 4412
rect 240 4222 2524 4256
rect 240 4066 2524 4100
rect 240 3910 2524 3944
rect 240 3754 2524 3788
rect 240 3598 2524 3632
rect 240 3442 2524 3476
rect 240 3286 2524 3320
rect 240 3130 2524 3164
rect 240 2974 2524 3008
rect 240 2818 2524 2852
rect 240 2662 2524 2696
rect 240 2506 2524 2540
rect 240 2350 2524 2384
rect 240 2194 2524 2228
rect 240 2038 2524 2072
rect 240 1882 2524 1916
rect 240 1726 2524 1760
rect 240 1570 2524 1604
rect 240 1414 2524 1448
rect 240 1258 2524 1292
rect 240 1102 2524 1136
rect 240 946 2524 980
rect 240 790 2524 824
rect 240 634 2524 668
rect 240 478 2524 512
rect 240 322 2524 356
rect 240 166 2524 200
<< mvnsubdiff >>
rect 66 43010 130 43044
rect 2556 43010 2620 43044
rect 66 42980 100 43010
rect 2586 42980 2620 43010
rect 66 100 100 130
rect 2586 100 2620 130
rect 66 66 130 100
rect 2556 66 2620 100
<< mvnsubdiffcont >>
rect 130 43010 2556 43044
rect 66 130 100 42980
rect 2586 130 2620 42980
rect 130 66 2556 100
<< poly >>
rect 140 42867 232 42899
rect 140 243 150 42867
rect 184 42799 232 42867
rect 2532 42799 2558 42899
rect 184 42743 217 42799
rect 184 42643 232 42743
rect 2532 42643 2558 42743
rect 184 42587 217 42643
rect 184 42487 232 42587
rect 2532 42487 2558 42587
rect 184 42431 217 42487
rect 184 42331 232 42431
rect 2532 42331 2558 42431
rect 184 42275 217 42331
rect 184 42175 232 42275
rect 2532 42175 2558 42275
rect 184 42119 217 42175
rect 184 42019 232 42119
rect 2532 42019 2558 42119
rect 184 41963 217 42019
rect 184 41863 232 41963
rect 2532 41863 2558 41963
rect 184 41807 217 41863
rect 184 41707 232 41807
rect 2532 41707 2558 41807
rect 184 41651 217 41707
rect 184 41551 232 41651
rect 2532 41551 2558 41651
rect 184 41495 217 41551
rect 184 41395 232 41495
rect 2532 41395 2558 41495
rect 184 41339 217 41395
rect 184 41239 232 41339
rect 2532 41239 2558 41339
rect 184 41183 217 41239
rect 184 41083 232 41183
rect 2532 41083 2558 41183
rect 184 41027 217 41083
rect 184 40927 232 41027
rect 2532 40927 2558 41027
rect 184 40871 217 40927
rect 184 40771 232 40871
rect 2532 40771 2558 40871
rect 184 40715 217 40771
rect 184 40615 232 40715
rect 2532 40615 2558 40715
rect 184 40559 217 40615
rect 184 40459 232 40559
rect 2532 40459 2558 40559
rect 184 40403 217 40459
rect 184 40303 232 40403
rect 2532 40303 2558 40403
rect 184 40247 217 40303
rect 184 40147 232 40247
rect 2532 40147 2558 40247
rect 184 40091 217 40147
rect 184 39991 232 40091
rect 2532 39991 2558 40091
rect 184 39935 217 39991
rect 184 39835 232 39935
rect 2532 39835 2558 39935
rect 184 39779 217 39835
rect 184 39679 232 39779
rect 2532 39679 2558 39779
rect 184 39623 217 39679
rect 184 39523 232 39623
rect 2532 39523 2558 39623
rect 184 39467 217 39523
rect 184 39367 232 39467
rect 2532 39367 2558 39467
rect 184 39311 217 39367
rect 184 39211 232 39311
rect 2532 39211 2558 39311
rect 184 39155 217 39211
rect 184 39055 232 39155
rect 2532 39055 2558 39155
rect 184 38999 217 39055
rect 184 38899 232 38999
rect 2532 38899 2558 38999
rect 184 38843 217 38899
rect 184 38743 232 38843
rect 2532 38743 2558 38843
rect 184 38687 217 38743
rect 184 38587 232 38687
rect 2532 38587 2558 38687
rect 184 38531 217 38587
rect 184 38431 232 38531
rect 2532 38431 2558 38531
rect 184 38375 217 38431
rect 184 38275 232 38375
rect 2532 38275 2558 38375
rect 184 38219 217 38275
rect 184 38119 232 38219
rect 2532 38119 2558 38219
rect 184 38063 217 38119
rect 184 37963 232 38063
rect 2532 37963 2558 38063
rect 184 37907 217 37963
rect 184 37807 232 37907
rect 2532 37807 2558 37907
rect 184 37751 217 37807
rect 184 37651 232 37751
rect 2532 37651 2558 37751
rect 184 37595 217 37651
rect 184 37495 232 37595
rect 2532 37495 2558 37595
rect 184 37439 217 37495
rect 184 37339 232 37439
rect 2532 37339 2558 37439
rect 184 37283 217 37339
rect 184 37183 232 37283
rect 2532 37183 2558 37283
rect 184 37127 217 37183
rect 184 37027 232 37127
rect 2532 37027 2558 37127
rect 184 36971 217 37027
rect 184 36871 232 36971
rect 2532 36871 2558 36971
rect 184 36815 217 36871
rect 184 36715 232 36815
rect 2532 36715 2558 36815
rect 184 36659 217 36715
rect 184 36559 232 36659
rect 2532 36559 2558 36659
rect 184 36503 217 36559
rect 184 36403 232 36503
rect 2532 36403 2558 36503
rect 184 36347 217 36403
rect 184 36247 232 36347
rect 2532 36247 2558 36347
rect 184 36191 217 36247
rect 184 36091 232 36191
rect 2532 36091 2558 36191
rect 184 36035 217 36091
rect 184 35935 232 36035
rect 2532 35935 2558 36035
rect 184 35879 217 35935
rect 184 35779 232 35879
rect 2532 35779 2558 35879
rect 184 35723 217 35779
rect 184 35623 232 35723
rect 2532 35623 2558 35723
rect 184 35567 217 35623
rect 184 35467 232 35567
rect 2532 35467 2558 35567
rect 184 35411 217 35467
rect 184 35311 232 35411
rect 2532 35311 2558 35411
rect 184 35255 217 35311
rect 184 35155 232 35255
rect 2532 35155 2558 35255
rect 184 35099 217 35155
rect 184 34999 232 35099
rect 2532 34999 2558 35099
rect 184 34943 217 34999
rect 184 34843 232 34943
rect 2532 34843 2558 34943
rect 184 34787 217 34843
rect 184 34687 232 34787
rect 2532 34687 2558 34787
rect 184 34631 217 34687
rect 184 34531 232 34631
rect 2532 34531 2558 34631
rect 184 34475 217 34531
rect 184 34375 232 34475
rect 2532 34375 2558 34475
rect 184 34319 217 34375
rect 184 34219 232 34319
rect 2532 34219 2558 34319
rect 184 34163 217 34219
rect 184 34063 232 34163
rect 2532 34063 2558 34163
rect 184 34007 217 34063
rect 184 33907 232 34007
rect 2532 33907 2558 34007
rect 184 33851 217 33907
rect 184 33751 232 33851
rect 2532 33751 2558 33851
rect 184 33695 217 33751
rect 184 33595 232 33695
rect 2532 33595 2558 33695
rect 184 33539 217 33595
rect 184 33439 232 33539
rect 2532 33439 2558 33539
rect 184 33383 217 33439
rect 184 33283 232 33383
rect 2532 33283 2558 33383
rect 184 33227 217 33283
rect 184 33127 232 33227
rect 2532 33127 2558 33227
rect 184 33071 217 33127
rect 184 32971 232 33071
rect 2532 32971 2558 33071
rect 184 32915 217 32971
rect 184 32815 232 32915
rect 2532 32815 2558 32915
rect 184 32759 217 32815
rect 184 32659 232 32759
rect 2532 32659 2558 32759
rect 184 32603 217 32659
rect 184 32503 232 32603
rect 2532 32503 2558 32603
rect 184 32447 217 32503
rect 184 32347 232 32447
rect 2532 32347 2558 32447
rect 184 32291 217 32347
rect 184 32191 232 32291
rect 2532 32191 2558 32291
rect 184 32135 217 32191
rect 184 32035 232 32135
rect 2532 32035 2558 32135
rect 184 31979 217 32035
rect 184 31879 232 31979
rect 2532 31879 2558 31979
rect 184 31823 217 31879
rect 184 31723 232 31823
rect 2532 31723 2558 31823
rect 184 31667 217 31723
rect 184 31567 232 31667
rect 2532 31567 2558 31667
rect 184 31511 217 31567
rect 184 31411 232 31511
rect 2532 31411 2558 31511
rect 184 31355 217 31411
rect 184 31255 232 31355
rect 2532 31255 2558 31355
rect 184 31199 217 31255
rect 184 31099 232 31199
rect 2532 31099 2558 31199
rect 184 31043 217 31099
rect 184 30943 232 31043
rect 2532 30943 2558 31043
rect 184 30887 217 30943
rect 184 30787 232 30887
rect 2532 30787 2558 30887
rect 184 30731 217 30787
rect 184 30631 232 30731
rect 2532 30631 2558 30731
rect 184 30575 217 30631
rect 184 30475 232 30575
rect 2532 30475 2558 30575
rect 184 30419 217 30475
rect 184 30319 232 30419
rect 2532 30319 2558 30419
rect 184 30263 217 30319
rect 184 30163 232 30263
rect 2532 30163 2558 30263
rect 184 30107 217 30163
rect 184 30007 232 30107
rect 2532 30007 2558 30107
rect 184 29951 217 30007
rect 184 29851 232 29951
rect 2532 29851 2558 29951
rect 184 29795 217 29851
rect 184 29695 232 29795
rect 2532 29695 2558 29795
rect 184 29639 217 29695
rect 184 29539 232 29639
rect 2532 29539 2558 29639
rect 184 29483 217 29539
rect 184 29383 232 29483
rect 2532 29383 2558 29483
rect 184 29327 217 29383
rect 184 29227 232 29327
rect 2532 29227 2558 29327
rect 184 29171 217 29227
rect 184 29071 232 29171
rect 2532 29071 2558 29171
rect 184 29015 217 29071
rect 184 28915 232 29015
rect 2532 28915 2558 29015
rect 184 28859 217 28915
rect 184 28759 232 28859
rect 2532 28759 2558 28859
rect 184 28703 217 28759
rect 184 28603 232 28703
rect 2532 28603 2558 28703
rect 184 28547 217 28603
rect 184 28447 232 28547
rect 2532 28447 2558 28547
rect 184 28391 217 28447
rect 184 28291 232 28391
rect 2532 28291 2558 28391
rect 184 28235 217 28291
rect 184 28135 232 28235
rect 2532 28135 2558 28235
rect 184 28079 217 28135
rect 184 27979 232 28079
rect 2532 27979 2558 28079
rect 184 27923 217 27979
rect 184 27823 232 27923
rect 2532 27823 2558 27923
rect 184 27767 217 27823
rect 184 27667 232 27767
rect 2532 27667 2558 27767
rect 184 27611 217 27667
rect 184 27511 232 27611
rect 2532 27511 2558 27611
rect 184 27455 217 27511
rect 184 27355 232 27455
rect 2532 27355 2558 27455
rect 184 27299 217 27355
rect 184 27199 232 27299
rect 2532 27199 2558 27299
rect 184 27143 217 27199
rect 184 27043 232 27143
rect 2532 27043 2558 27143
rect 184 26987 217 27043
rect 184 26887 232 26987
rect 2532 26887 2558 26987
rect 184 26831 217 26887
rect 184 26731 232 26831
rect 2532 26731 2558 26831
rect 184 26675 217 26731
rect 184 26575 232 26675
rect 2532 26575 2558 26675
rect 184 26519 217 26575
rect 184 26419 232 26519
rect 2532 26419 2558 26519
rect 184 26363 217 26419
rect 184 26263 232 26363
rect 2532 26263 2558 26363
rect 184 26207 217 26263
rect 184 26107 232 26207
rect 2532 26107 2558 26207
rect 184 26051 217 26107
rect 184 25951 232 26051
rect 2532 25951 2558 26051
rect 184 25895 217 25951
rect 184 25795 232 25895
rect 2532 25795 2558 25895
rect 184 25739 217 25795
rect 184 25639 232 25739
rect 2532 25639 2558 25739
rect 184 25583 217 25639
rect 184 25483 232 25583
rect 2532 25483 2558 25583
rect 184 25427 217 25483
rect 184 25327 232 25427
rect 2532 25327 2558 25427
rect 184 25271 217 25327
rect 184 25171 232 25271
rect 2532 25171 2558 25271
rect 184 25115 217 25171
rect 184 25015 232 25115
rect 2532 25015 2558 25115
rect 184 24959 217 25015
rect 184 24859 232 24959
rect 2532 24859 2558 24959
rect 184 24803 217 24859
rect 184 24703 232 24803
rect 2532 24703 2558 24803
rect 184 24647 217 24703
rect 184 24547 232 24647
rect 2532 24547 2558 24647
rect 184 24491 217 24547
rect 184 24391 232 24491
rect 2532 24391 2558 24491
rect 184 24335 217 24391
rect 184 24235 232 24335
rect 2532 24235 2558 24335
rect 184 24179 217 24235
rect 184 24079 232 24179
rect 2532 24079 2558 24179
rect 184 24023 217 24079
rect 184 23923 232 24023
rect 2532 23923 2558 24023
rect 184 23867 217 23923
rect 184 23767 232 23867
rect 2532 23767 2558 23867
rect 184 23711 217 23767
rect 184 23611 232 23711
rect 2532 23611 2558 23711
rect 184 23555 217 23611
rect 184 23455 232 23555
rect 2532 23455 2558 23555
rect 184 23399 217 23455
rect 184 23299 232 23399
rect 2532 23299 2558 23399
rect 184 23243 217 23299
rect 184 23143 232 23243
rect 2532 23143 2558 23243
rect 184 23087 217 23143
rect 184 22987 232 23087
rect 2532 22987 2558 23087
rect 184 22931 217 22987
rect 184 22831 232 22931
rect 2532 22831 2558 22931
rect 184 22775 217 22831
rect 184 22675 232 22775
rect 2532 22675 2558 22775
rect 184 22619 217 22675
rect 184 22519 232 22619
rect 2532 22519 2558 22619
rect 184 22463 217 22519
rect 184 22363 232 22463
rect 2532 22363 2558 22463
rect 184 22307 217 22363
rect 184 22207 232 22307
rect 2532 22207 2558 22307
rect 184 22151 217 22207
rect 184 22051 232 22151
rect 2532 22051 2558 22151
rect 184 21995 217 22051
rect 184 21895 232 21995
rect 2532 21895 2558 21995
rect 184 21839 217 21895
rect 184 21739 232 21839
rect 2532 21739 2558 21839
rect 184 21683 217 21739
rect 184 21583 232 21683
rect 2532 21583 2558 21683
rect 184 21527 217 21583
rect 184 21427 232 21527
rect 2532 21427 2558 21527
rect 184 21371 217 21427
rect 184 21271 232 21371
rect 2532 21271 2558 21371
rect 184 21215 217 21271
rect 184 21115 232 21215
rect 2532 21115 2558 21215
rect 184 21059 217 21115
rect 184 20959 232 21059
rect 2532 20959 2558 21059
rect 184 20903 217 20959
rect 184 20803 232 20903
rect 2532 20803 2558 20903
rect 184 20747 217 20803
rect 184 20647 232 20747
rect 2532 20647 2558 20747
rect 184 20591 217 20647
rect 184 20491 232 20591
rect 2532 20491 2558 20591
rect 184 20435 217 20491
rect 184 20335 232 20435
rect 2532 20335 2558 20435
rect 184 20279 217 20335
rect 184 20179 232 20279
rect 2532 20179 2558 20279
rect 184 20123 217 20179
rect 184 20023 232 20123
rect 2532 20023 2558 20123
rect 184 19967 217 20023
rect 184 19867 232 19967
rect 2532 19867 2558 19967
rect 184 19811 217 19867
rect 184 19711 232 19811
rect 2532 19711 2558 19811
rect 184 19655 217 19711
rect 184 19555 232 19655
rect 2532 19555 2558 19655
rect 184 19499 217 19555
rect 184 19399 232 19499
rect 2532 19399 2558 19499
rect 184 19343 217 19399
rect 184 19243 232 19343
rect 2532 19243 2558 19343
rect 184 19187 217 19243
rect 184 19087 232 19187
rect 2532 19087 2558 19187
rect 184 19031 217 19087
rect 184 18931 232 19031
rect 2532 18931 2558 19031
rect 184 18875 217 18931
rect 184 18775 232 18875
rect 2532 18775 2558 18875
rect 184 18719 217 18775
rect 184 18619 232 18719
rect 2532 18619 2558 18719
rect 184 18563 217 18619
rect 184 18463 232 18563
rect 2532 18463 2558 18563
rect 184 18407 217 18463
rect 184 18307 232 18407
rect 2532 18307 2558 18407
rect 184 18251 217 18307
rect 184 18151 232 18251
rect 2532 18151 2558 18251
rect 184 18095 217 18151
rect 184 17995 232 18095
rect 2532 17995 2558 18095
rect 184 17939 217 17995
rect 184 17839 232 17939
rect 2532 17839 2558 17939
rect 184 17783 217 17839
rect 184 17683 232 17783
rect 2532 17683 2558 17783
rect 184 17627 217 17683
rect 184 17527 232 17627
rect 2532 17527 2558 17627
rect 184 17471 217 17527
rect 184 17371 232 17471
rect 2532 17371 2558 17471
rect 184 17315 217 17371
rect 184 17215 232 17315
rect 2532 17215 2558 17315
rect 184 17159 217 17215
rect 184 17059 232 17159
rect 2532 17059 2558 17159
rect 184 17003 217 17059
rect 184 16903 232 17003
rect 2532 16903 2558 17003
rect 184 16847 217 16903
rect 184 16747 232 16847
rect 2532 16747 2558 16847
rect 184 16691 217 16747
rect 184 16591 232 16691
rect 2532 16591 2558 16691
rect 184 16535 217 16591
rect 184 16435 232 16535
rect 2532 16435 2558 16535
rect 184 16379 217 16435
rect 184 16279 232 16379
rect 2532 16279 2558 16379
rect 184 16223 217 16279
rect 184 16123 232 16223
rect 2532 16123 2558 16223
rect 184 16067 217 16123
rect 184 15967 232 16067
rect 2532 15967 2558 16067
rect 184 15911 217 15967
rect 184 15811 232 15911
rect 2532 15811 2558 15911
rect 184 15755 217 15811
rect 184 15655 232 15755
rect 2532 15655 2558 15755
rect 184 15599 217 15655
rect 184 15499 232 15599
rect 2532 15499 2558 15599
rect 184 15443 217 15499
rect 184 15343 232 15443
rect 2532 15343 2558 15443
rect 184 15287 217 15343
rect 184 15187 232 15287
rect 2532 15187 2558 15287
rect 184 15131 217 15187
rect 184 15031 232 15131
rect 2532 15031 2558 15131
rect 184 14975 217 15031
rect 184 14875 232 14975
rect 2532 14875 2558 14975
rect 184 14819 217 14875
rect 184 14719 232 14819
rect 2532 14719 2558 14819
rect 184 14663 217 14719
rect 184 14563 232 14663
rect 2532 14563 2558 14663
rect 184 14507 217 14563
rect 184 14407 232 14507
rect 2532 14407 2558 14507
rect 184 14351 217 14407
rect 184 14251 232 14351
rect 2532 14251 2558 14351
rect 184 14195 217 14251
rect 184 14095 232 14195
rect 2532 14095 2558 14195
rect 184 14039 217 14095
rect 184 13939 232 14039
rect 2532 13939 2558 14039
rect 184 13883 217 13939
rect 184 13783 232 13883
rect 2532 13783 2558 13883
rect 184 13727 217 13783
rect 184 13627 232 13727
rect 2532 13627 2558 13727
rect 184 13571 217 13627
rect 184 13471 232 13571
rect 2532 13471 2558 13571
rect 184 13415 217 13471
rect 184 13315 232 13415
rect 2532 13315 2558 13415
rect 184 13259 217 13315
rect 184 13159 232 13259
rect 2532 13159 2558 13259
rect 184 13103 217 13159
rect 184 13003 232 13103
rect 2532 13003 2558 13103
rect 184 12947 217 13003
rect 184 12847 232 12947
rect 2532 12847 2558 12947
rect 184 12791 217 12847
rect 184 12691 232 12791
rect 2532 12691 2558 12791
rect 184 12635 217 12691
rect 184 12535 232 12635
rect 2532 12535 2558 12635
rect 184 12479 217 12535
rect 184 12379 232 12479
rect 2532 12379 2558 12479
rect 184 12323 217 12379
rect 184 12223 232 12323
rect 2532 12223 2558 12323
rect 184 12167 217 12223
rect 184 12067 232 12167
rect 2532 12067 2558 12167
rect 184 12011 217 12067
rect 184 11911 232 12011
rect 2532 11911 2558 12011
rect 184 11855 217 11911
rect 184 11755 232 11855
rect 2532 11755 2558 11855
rect 184 11699 217 11755
rect 184 11599 232 11699
rect 2532 11599 2558 11699
rect 184 11543 217 11599
rect 184 11443 232 11543
rect 2532 11443 2558 11543
rect 184 11387 217 11443
rect 184 11287 232 11387
rect 2532 11287 2558 11387
rect 184 11231 217 11287
rect 184 11131 232 11231
rect 2532 11131 2558 11231
rect 184 11075 217 11131
rect 184 10975 232 11075
rect 2532 10975 2558 11075
rect 184 10919 217 10975
rect 184 10819 232 10919
rect 2532 10819 2558 10919
rect 184 10763 217 10819
rect 184 10663 232 10763
rect 2532 10663 2558 10763
rect 184 10607 217 10663
rect 184 10507 232 10607
rect 2532 10507 2558 10607
rect 184 10451 217 10507
rect 184 10351 232 10451
rect 2532 10351 2558 10451
rect 184 10295 217 10351
rect 184 10195 232 10295
rect 2532 10195 2558 10295
rect 184 10139 217 10195
rect 184 10039 232 10139
rect 2532 10039 2558 10139
rect 184 9983 217 10039
rect 184 9883 232 9983
rect 2532 9883 2558 9983
rect 184 9827 217 9883
rect 184 9727 232 9827
rect 2532 9727 2558 9827
rect 184 9671 217 9727
rect 184 9571 232 9671
rect 2532 9571 2558 9671
rect 184 9515 217 9571
rect 184 9415 232 9515
rect 2532 9415 2558 9515
rect 184 9359 217 9415
rect 184 9259 232 9359
rect 2532 9259 2558 9359
rect 184 9203 217 9259
rect 184 9103 232 9203
rect 2532 9103 2558 9203
rect 184 9047 217 9103
rect 184 8947 232 9047
rect 2532 8947 2558 9047
rect 184 8891 217 8947
rect 184 8791 232 8891
rect 2532 8791 2558 8891
rect 184 8735 217 8791
rect 184 8635 232 8735
rect 2532 8635 2558 8735
rect 184 8579 217 8635
rect 184 8479 232 8579
rect 2532 8479 2558 8579
rect 184 8423 217 8479
rect 184 8323 232 8423
rect 2532 8323 2558 8423
rect 184 8267 217 8323
rect 184 8167 232 8267
rect 2532 8167 2558 8267
rect 184 8111 217 8167
rect 184 8011 232 8111
rect 2532 8011 2558 8111
rect 184 7955 217 8011
rect 184 7855 232 7955
rect 2532 7855 2558 7955
rect 184 7799 217 7855
rect 184 7699 232 7799
rect 2532 7699 2558 7799
rect 184 7643 217 7699
rect 184 7543 232 7643
rect 2532 7543 2558 7643
rect 184 7487 217 7543
rect 184 7387 232 7487
rect 2532 7387 2558 7487
rect 184 7331 217 7387
rect 184 7231 232 7331
rect 2532 7231 2558 7331
rect 184 7175 217 7231
rect 184 7075 232 7175
rect 2532 7075 2558 7175
rect 184 7019 217 7075
rect 184 6919 232 7019
rect 2532 6919 2558 7019
rect 184 6863 217 6919
rect 184 6763 232 6863
rect 2532 6763 2558 6863
rect 184 6707 217 6763
rect 184 6607 232 6707
rect 2532 6607 2558 6707
rect 184 6551 217 6607
rect 184 6451 232 6551
rect 2532 6451 2558 6551
rect 184 6395 217 6451
rect 184 6295 232 6395
rect 2532 6295 2558 6395
rect 184 6239 217 6295
rect 184 6139 232 6239
rect 2532 6139 2558 6239
rect 184 6083 217 6139
rect 184 5983 232 6083
rect 2532 5983 2558 6083
rect 184 5927 217 5983
rect 184 5827 232 5927
rect 2532 5827 2558 5927
rect 184 5771 217 5827
rect 184 5671 232 5771
rect 2532 5671 2558 5771
rect 184 5615 217 5671
rect 184 5515 232 5615
rect 2532 5515 2558 5615
rect 184 5459 217 5515
rect 184 5359 232 5459
rect 2532 5359 2558 5459
rect 184 5303 217 5359
rect 184 5203 232 5303
rect 2532 5203 2558 5303
rect 184 5147 217 5203
rect 184 5047 232 5147
rect 2532 5047 2558 5147
rect 184 4991 217 5047
rect 184 4891 232 4991
rect 2532 4891 2558 4991
rect 184 4835 217 4891
rect 184 4735 232 4835
rect 2532 4735 2558 4835
rect 184 4679 217 4735
rect 184 4579 232 4679
rect 2532 4579 2558 4679
rect 184 4523 217 4579
rect 184 4423 232 4523
rect 2532 4423 2558 4523
rect 184 4367 217 4423
rect 184 4267 232 4367
rect 2532 4267 2558 4367
rect 184 4211 217 4267
rect 184 4111 232 4211
rect 2532 4111 2558 4211
rect 184 4055 217 4111
rect 184 3955 232 4055
rect 2532 3955 2558 4055
rect 184 3899 217 3955
rect 184 3799 232 3899
rect 2532 3799 2558 3899
rect 184 3743 217 3799
rect 184 3643 232 3743
rect 2532 3643 2558 3743
rect 184 3587 217 3643
rect 184 3487 232 3587
rect 2532 3487 2558 3587
rect 184 3431 217 3487
rect 184 3331 232 3431
rect 2532 3331 2558 3431
rect 184 3275 217 3331
rect 184 3175 232 3275
rect 2532 3175 2558 3275
rect 184 3119 217 3175
rect 184 3019 232 3119
rect 2532 3019 2558 3119
rect 184 2963 217 3019
rect 184 2863 232 2963
rect 2532 2863 2558 2963
rect 184 2807 217 2863
rect 184 2707 232 2807
rect 2532 2707 2558 2807
rect 184 2651 217 2707
rect 184 2551 232 2651
rect 2532 2551 2558 2651
rect 184 2495 217 2551
rect 184 2395 232 2495
rect 2532 2395 2558 2495
rect 184 2339 217 2395
rect 184 2239 232 2339
rect 2532 2239 2558 2339
rect 184 2183 217 2239
rect 184 2083 232 2183
rect 2532 2083 2558 2183
rect 184 2027 217 2083
rect 184 1927 232 2027
rect 2532 1927 2558 2027
rect 184 1871 217 1927
rect 184 1771 232 1871
rect 2532 1771 2558 1871
rect 184 1715 217 1771
rect 184 1615 232 1715
rect 2532 1615 2558 1715
rect 184 1559 217 1615
rect 184 1459 232 1559
rect 2532 1459 2558 1559
rect 184 1403 217 1459
rect 184 1303 232 1403
rect 2532 1303 2558 1403
rect 184 1247 217 1303
rect 184 1147 232 1247
rect 2532 1147 2558 1247
rect 184 1091 217 1147
rect 184 991 232 1091
rect 2532 991 2558 1091
rect 184 935 217 991
rect 184 835 232 935
rect 2532 835 2558 935
rect 184 779 217 835
rect 184 679 232 779
rect 2532 679 2558 779
rect 184 623 217 679
rect 184 523 232 623
rect 2532 523 2558 623
rect 184 467 217 523
rect 184 367 232 467
rect 2532 367 2558 467
rect 184 311 217 367
rect 184 243 232 311
rect 140 211 232 243
rect 2532 211 2558 311
<< polycont >>
rect 150 243 184 42867
<< locali >>
rect 66 43010 130 43044
rect 2556 43010 2620 43044
rect 66 42980 100 43010
rect 2586 42980 2620 43010
rect 224 42910 240 42944
rect 2524 42910 2540 42944
rect 150 42871 184 42883
rect 224 42754 240 42788
rect 2524 42754 2540 42788
rect 224 42598 240 42632
rect 2524 42598 2540 42632
rect 224 42442 240 42476
rect 2524 42442 2540 42476
rect 224 42286 240 42320
rect 2524 42286 2540 42320
rect 224 42130 240 42164
rect 2524 42130 2540 42164
rect 224 41974 240 42008
rect 2524 41974 2540 42008
rect 224 41818 240 41852
rect 2524 41818 2540 41852
rect 224 41662 240 41696
rect 2524 41662 2540 41696
rect 224 41506 240 41540
rect 2524 41506 2540 41540
rect 224 41350 240 41384
rect 2524 41350 2540 41384
rect 224 41194 240 41228
rect 2524 41194 2540 41228
rect 224 41038 240 41072
rect 2524 41038 2540 41072
rect 224 40882 240 40916
rect 2524 40882 2540 40916
rect 224 40726 240 40760
rect 2524 40726 2540 40760
rect 224 40570 240 40604
rect 2524 40570 2540 40604
rect 224 40414 240 40448
rect 2524 40414 2540 40448
rect 224 40258 240 40292
rect 2524 40258 2540 40292
rect 224 40102 240 40136
rect 2524 40102 2540 40136
rect 224 39946 240 39980
rect 2524 39946 2540 39980
rect 224 39790 240 39824
rect 2524 39790 2540 39824
rect 224 39634 240 39668
rect 2524 39634 2540 39668
rect 224 39478 240 39512
rect 2524 39478 2540 39512
rect 224 39322 240 39356
rect 2524 39322 2540 39356
rect 224 39166 240 39200
rect 2524 39166 2540 39200
rect 224 39010 240 39044
rect 2524 39010 2540 39044
rect 224 38854 240 38888
rect 2524 38854 2540 38888
rect 224 38698 240 38732
rect 2524 38698 2540 38732
rect 224 38542 240 38576
rect 2524 38542 2540 38576
rect 224 38386 240 38420
rect 2524 38386 2540 38420
rect 224 38230 240 38264
rect 2524 38230 2540 38264
rect 224 38074 240 38108
rect 2524 38074 2540 38108
rect 224 37918 240 37952
rect 2524 37918 2540 37952
rect 224 37762 240 37796
rect 2524 37762 2540 37796
rect 224 37606 240 37640
rect 2524 37606 2540 37640
rect 224 37450 240 37484
rect 2524 37450 2540 37484
rect 224 37294 240 37328
rect 2524 37294 2540 37328
rect 224 37138 240 37172
rect 2524 37138 2540 37172
rect 224 36982 240 37016
rect 2524 36982 2540 37016
rect 224 36826 240 36860
rect 2524 36826 2540 36860
rect 224 36670 240 36704
rect 2524 36670 2540 36704
rect 224 36514 240 36548
rect 2524 36514 2540 36548
rect 224 36358 240 36392
rect 2524 36358 2540 36392
rect 224 36202 240 36236
rect 2524 36202 2540 36236
rect 224 36046 240 36080
rect 2524 36046 2540 36080
rect 224 35890 240 35924
rect 2524 35890 2540 35924
rect 224 35734 240 35768
rect 2524 35734 2540 35768
rect 224 35578 240 35612
rect 2524 35578 2540 35612
rect 224 35422 240 35456
rect 2524 35422 2540 35456
rect 224 35266 240 35300
rect 2524 35266 2540 35300
rect 224 35110 240 35144
rect 2524 35110 2540 35144
rect 224 34954 240 34988
rect 2524 34954 2540 34988
rect 224 34798 240 34832
rect 2524 34798 2540 34832
rect 224 34642 240 34676
rect 2524 34642 2540 34676
rect 224 34486 240 34520
rect 2524 34486 2540 34520
rect 224 34330 240 34364
rect 2524 34330 2540 34364
rect 224 34174 240 34208
rect 2524 34174 2540 34208
rect 224 34018 240 34052
rect 2524 34018 2540 34052
rect 224 33862 240 33896
rect 2524 33862 2540 33896
rect 224 33706 240 33740
rect 2524 33706 2540 33740
rect 224 33550 240 33584
rect 2524 33550 2540 33584
rect 224 33394 240 33428
rect 2524 33394 2540 33428
rect 224 33238 240 33272
rect 2524 33238 2540 33272
rect 224 33082 240 33116
rect 2524 33082 2540 33116
rect 224 32926 240 32960
rect 2524 32926 2540 32960
rect 224 32770 240 32804
rect 2524 32770 2540 32804
rect 224 32614 240 32648
rect 2524 32614 2540 32648
rect 224 32458 240 32492
rect 2524 32458 2540 32492
rect 224 32302 240 32336
rect 2524 32302 2540 32336
rect 224 32146 240 32180
rect 2524 32146 2540 32180
rect 224 31990 240 32024
rect 2524 31990 2540 32024
rect 224 31834 240 31868
rect 2524 31834 2540 31868
rect 224 31678 240 31712
rect 2524 31678 2540 31712
rect 224 31522 240 31556
rect 2524 31522 2540 31556
rect 224 31366 240 31400
rect 2524 31366 2540 31400
rect 224 31210 240 31244
rect 2524 31210 2540 31244
rect 224 31054 240 31088
rect 2524 31054 2540 31088
rect 224 30898 240 30932
rect 2524 30898 2540 30932
rect 224 30742 240 30776
rect 2524 30742 2540 30776
rect 224 30586 240 30620
rect 2524 30586 2540 30620
rect 224 30430 240 30464
rect 2524 30430 2540 30464
rect 224 30274 240 30308
rect 2524 30274 2540 30308
rect 224 30118 240 30152
rect 2524 30118 2540 30152
rect 224 29962 240 29996
rect 2524 29962 2540 29996
rect 224 29806 240 29840
rect 2524 29806 2540 29840
rect 224 29650 240 29684
rect 2524 29650 2540 29684
rect 224 29494 240 29528
rect 2524 29494 2540 29528
rect 224 29338 240 29372
rect 2524 29338 2540 29372
rect 224 29182 240 29216
rect 2524 29182 2540 29216
rect 224 29026 240 29060
rect 2524 29026 2540 29060
rect 224 28870 240 28904
rect 2524 28870 2540 28904
rect 224 28714 240 28748
rect 2524 28714 2540 28748
rect 224 28558 240 28592
rect 2524 28558 2540 28592
rect 224 28402 240 28436
rect 2524 28402 2540 28436
rect 224 28246 240 28280
rect 2524 28246 2540 28280
rect 224 28090 240 28124
rect 2524 28090 2540 28124
rect 224 27934 240 27968
rect 2524 27934 2540 27968
rect 224 27778 240 27812
rect 2524 27778 2540 27812
rect 224 27622 240 27656
rect 2524 27622 2540 27656
rect 224 27466 240 27500
rect 2524 27466 2540 27500
rect 224 27310 240 27344
rect 2524 27310 2540 27344
rect 224 27154 240 27188
rect 2524 27154 2540 27188
rect 224 26998 240 27032
rect 2524 26998 2540 27032
rect 224 26842 240 26876
rect 2524 26842 2540 26876
rect 224 26686 240 26720
rect 2524 26686 2540 26720
rect 224 26530 240 26564
rect 2524 26530 2540 26564
rect 224 26374 240 26408
rect 2524 26374 2540 26408
rect 224 26218 240 26252
rect 2524 26218 2540 26252
rect 224 26062 240 26096
rect 2524 26062 2540 26096
rect 224 25906 240 25940
rect 2524 25906 2540 25940
rect 224 25750 240 25784
rect 2524 25750 2540 25784
rect 224 25594 240 25628
rect 2524 25594 2540 25628
rect 224 25438 240 25472
rect 2524 25438 2540 25472
rect 224 25282 240 25316
rect 2524 25282 2540 25316
rect 224 25126 240 25160
rect 2524 25126 2540 25160
rect 224 24970 240 25004
rect 2524 24970 2540 25004
rect 224 24814 240 24848
rect 2524 24814 2540 24848
rect 224 24658 240 24692
rect 2524 24658 2540 24692
rect 224 24502 240 24536
rect 2524 24502 2540 24536
rect 224 24346 240 24380
rect 2524 24346 2540 24380
rect 224 24190 240 24224
rect 2524 24190 2540 24224
rect 224 24034 240 24068
rect 2524 24034 2540 24068
rect 224 23878 240 23912
rect 2524 23878 2540 23912
rect 224 23722 240 23756
rect 2524 23722 2540 23756
rect 224 23566 240 23600
rect 2524 23566 2540 23600
rect 224 23410 240 23444
rect 2524 23410 2540 23444
rect 224 23254 240 23288
rect 2524 23254 2540 23288
rect 224 23098 240 23132
rect 2524 23098 2540 23132
rect 224 22942 240 22976
rect 2524 22942 2540 22976
rect 224 22786 240 22820
rect 2524 22786 2540 22820
rect 224 22630 240 22664
rect 2524 22630 2540 22664
rect 224 22474 240 22508
rect 2524 22474 2540 22508
rect 224 22318 240 22352
rect 2524 22318 2540 22352
rect 224 22162 240 22196
rect 2524 22162 2540 22196
rect 224 22006 240 22040
rect 2524 22006 2540 22040
rect 224 21850 240 21884
rect 2524 21850 2540 21884
rect 224 21694 240 21728
rect 2524 21694 2540 21728
rect 224 21538 240 21572
rect 2524 21538 2540 21572
rect 224 21382 240 21416
rect 2524 21382 2540 21416
rect 224 21226 240 21260
rect 2524 21226 2540 21260
rect 224 21070 240 21104
rect 2524 21070 2540 21104
rect 224 20914 240 20948
rect 2524 20914 2540 20948
rect 224 20758 240 20792
rect 2524 20758 2540 20792
rect 224 20602 240 20636
rect 2524 20602 2540 20636
rect 224 20446 240 20480
rect 2524 20446 2540 20480
rect 224 20290 240 20324
rect 2524 20290 2540 20324
rect 224 20134 240 20168
rect 2524 20134 2540 20168
rect 224 19978 240 20012
rect 2524 19978 2540 20012
rect 224 19822 240 19856
rect 2524 19822 2540 19856
rect 224 19666 240 19700
rect 2524 19666 2540 19700
rect 224 19510 240 19544
rect 2524 19510 2540 19544
rect 224 19354 240 19388
rect 2524 19354 2540 19388
rect 224 19198 240 19232
rect 2524 19198 2540 19232
rect 224 19042 240 19076
rect 2524 19042 2540 19076
rect 224 18886 240 18920
rect 2524 18886 2540 18920
rect 224 18730 240 18764
rect 2524 18730 2540 18764
rect 224 18574 240 18608
rect 2524 18574 2540 18608
rect 224 18418 240 18452
rect 2524 18418 2540 18452
rect 224 18262 240 18296
rect 2524 18262 2540 18296
rect 224 18106 240 18140
rect 2524 18106 2540 18140
rect 224 17950 240 17984
rect 2524 17950 2540 17984
rect 224 17794 240 17828
rect 2524 17794 2540 17828
rect 224 17638 240 17672
rect 2524 17638 2540 17672
rect 224 17482 240 17516
rect 2524 17482 2540 17516
rect 224 17326 240 17360
rect 2524 17326 2540 17360
rect 224 17170 240 17204
rect 2524 17170 2540 17204
rect 224 17014 240 17048
rect 2524 17014 2540 17048
rect 224 16858 240 16892
rect 2524 16858 2540 16892
rect 224 16702 240 16736
rect 2524 16702 2540 16736
rect 224 16546 240 16580
rect 2524 16546 2540 16580
rect 224 16390 240 16424
rect 2524 16390 2540 16424
rect 224 16234 240 16268
rect 2524 16234 2540 16268
rect 224 16078 240 16112
rect 2524 16078 2540 16112
rect 224 15922 240 15956
rect 2524 15922 2540 15956
rect 224 15766 240 15800
rect 2524 15766 2540 15800
rect 224 15610 240 15644
rect 2524 15610 2540 15644
rect 224 15454 240 15488
rect 2524 15454 2540 15488
rect 224 15298 240 15332
rect 2524 15298 2540 15332
rect 224 15142 240 15176
rect 2524 15142 2540 15176
rect 224 14986 240 15020
rect 2524 14986 2540 15020
rect 224 14830 240 14864
rect 2524 14830 2540 14864
rect 224 14674 240 14708
rect 2524 14674 2540 14708
rect 224 14518 240 14552
rect 2524 14518 2540 14552
rect 224 14362 240 14396
rect 2524 14362 2540 14396
rect 224 14206 240 14240
rect 2524 14206 2540 14240
rect 224 14050 240 14084
rect 2524 14050 2540 14084
rect 224 13894 240 13928
rect 2524 13894 2540 13928
rect 224 13738 240 13772
rect 2524 13738 2540 13772
rect 224 13582 240 13616
rect 2524 13582 2540 13616
rect 224 13426 240 13460
rect 2524 13426 2540 13460
rect 224 13270 240 13304
rect 2524 13270 2540 13304
rect 224 13114 240 13148
rect 2524 13114 2540 13148
rect 224 12958 240 12992
rect 2524 12958 2540 12992
rect 224 12802 240 12836
rect 2524 12802 2540 12836
rect 224 12646 240 12680
rect 2524 12646 2540 12680
rect 224 12490 240 12524
rect 2524 12490 2540 12524
rect 224 12334 240 12368
rect 2524 12334 2540 12368
rect 224 12178 240 12212
rect 2524 12178 2540 12212
rect 224 12022 240 12056
rect 2524 12022 2540 12056
rect 224 11866 240 11900
rect 2524 11866 2540 11900
rect 224 11710 240 11744
rect 2524 11710 2540 11744
rect 224 11554 240 11588
rect 2524 11554 2540 11588
rect 224 11398 240 11432
rect 2524 11398 2540 11432
rect 224 11242 240 11276
rect 2524 11242 2540 11276
rect 224 11086 240 11120
rect 2524 11086 2540 11120
rect 224 10930 240 10964
rect 2524 10930 2540 10964
rect 224 10774 240 10808
rect 2524 10774 2540 10808
rect 224 10618 240 10652
rect 2524 10618 2540 10652
rect 224 10462 240 10496
rect 2524 10462 2540 10496
rect 224 10306 240 10340
rect 2524 10306 2540 10340
rect 224 10150 240 10184
rect 2524 10150 2540 10184
rect 224 9994 240 10028
rect 2524 9994 2540 10028
rect 224 9838 240 9872
rect 2524 9838 2540 9872
rect 224 9682 240 9716
rect 2524 9682 2540 9716
rect 224 9526 240 9560
rect 2524 9526 2540 9560
rect 224 9370 240 9404
rect 2524 9370 2540 9404
rect 224 9214 240 9248
rect 2524 9214 2540 9248
rect 224 9058 240 9092
rect 2524 9058 2540 9092
rect 224 8902 240 8936
rect 2524 8902 2540 8936
rect 224 8746 240 8780
rect 2524 8746 2540 8780
rect 224 8590 240 8624
rect 2524 8590 2540 8624
rect 224 8434 240 8468
rect 2524 8434 2540 8468
rect 224 8278 240 8312
rect 2524 8278 2540 8312
rect 224 8122 240 8156
rect 2524 8122 2540 8156
rect 224 7966 240 8000
rect 2524 7966 2540 8000
rect 224 7810 240 7844
rect 2524 7810 2540 7844
rect 224 7654 240 7688
rect 2524 7654 2540 7688
rect 224 7498 240 7532
rect 2524 7498 2540 7532
rect 224 7342 240 7376
rect 2524 7342 2540 7376
rect 224 7186 240 7220
rect 2524 7186 2540 7220
rect 224 7030 240 7064
rect 2524 7030 2540 7064
rect 224 6874 240 6908
rect 2524 6874 2540 6908
rect 224 6718 240 6752
rect 2524 6718 2540 6752
rect 224 6562 240 6596
rect 2524 6562 2540 6596
rect 224 6406 240 6440
rect 2524 6406 2540 6440
rect 224 6250 240 6284
rect 2524 6250 2540 6284
rect 224 6094 240 6128
rect 2524 6094 2540 6128
rect 224 5938 240 5972
rect 2524 5938 2540 5972
rect 224 5782 240 5816
rect 2524 5782 2540 5816
rect 224 5626 240 5660
rect 2524 5626 2540 5660
rect 224 5470 240 5504
rect 2524 5470 2540 5504
rect 224 5314 240 5348
rect 2524 5314 2540 5348
rect 224 5158 240 5192
rect 2524 5158 2540 5192
rect 224 5002 240 5036
rect 2524 5002 2540 5036
rect 224 4846 240 4880
rect 2524 4846 2540 4880
rect 224 4690 240 4724
rect 2524 4690 2540 4724
rect 224 4534 240 4568
rect 2524 4534 2540 4568
rect 224 4378 240 4412
rect 2524 4378 2540 4412
rect 224 4222 240 4256
rect 2524 4222 2540 4256
rect 224 4066 240 4100
rect 2524 4066 2540 4100
rect 224 3910 240 3944
rect 2524 3910 2540 3944
rect 224 3754 240 3788
rect 2524 3754 2540 3788
rect 224 3598 240 3632
rect 2524 3598 2540 3632
rect 224 3442 240 3476
rect 2524 3442 2540 3476
rect 224 3286 240 3320
rect 2524 3286 2540 3320
rect 224 3130 240 3164
rect 2524 3130 2540 3164
rect 224 2974 240 3008
rect 2524 2974 2540 3008
rect 224 2818 240 2852
rect 2524 2818 2540 2852
rect 224 2662 240 2696
rect 2524 2662 2540 2696
rect 224 2506 240 2540
rect 2524 2506 2540 2540
rect 224 2350 240 2384
rect 2524 2350 2540 2384
rect 224 2194 240 2228
rect 2524 2194 2540 2228
rect 224 2038 240 2072
rect 2524 2038 2540 2072
rect 224 1882 240 1916
rect 2524 1882 2540 1916
rect 224 1726 240 1760
rect 2524 1726 2540 1760
rect 224 1570 240 1604
rect 2524 1570 2540 1604
rect 224 1414 240 1448
rect 2524 1414 2540 1448
rect 224 1258 240 1292
rect 2524 1258 2540 1292
rect 224 1102 240 1136
rect 2524 1102 2540 1136
rect 224 946 240 980
rect 2524 946 2540 980
rect 224 790 240 824
rect 2524 790 2540 824
rect 224 634 240 668
rect 2524 634 2540 668
rect 224 478 240 512
rect 2524 478 2540 512
rect 224 322 240 356
rect 2524 322 2540 356
rect 150 227 184 239
rect 224 166 240 200
rect 2524 166 2540 200
rect 66 100 100 130
rect 2586 100 2620 130
rect 66 66 130 100
rect 2556 66 2620 100
<< viali >>
rect 130 43010 2556 43044
rect 66 130 100 42980
rect 240 42910 2524 42944
rect 150 42867 184 42871
rect 150 243 184 42867
rect 240 42754 2524 42788
rect 240 42598 2524 42632
rect 240 42442 2524 42476
rect 240 42286 2524 42320
rect 240 42130 2524 42164
rect 240 41974 2524 42008
rect 240 41818 2524 41852
rect 240 41662 2524 41696
rect 240 41506 2524 41540
rect 240 41350 2524 41384
rect 240 41194 2524 41228
rect 240 41038 2524 41072
rect 240 40882 2524 40916
rect 240 40726 2524 40760
rect 240 40570 2524 40604
rect 240 40414 2524 40448
rect 240 40258 2524 40292
rect 240 40102 2524 40136
rect 240 39946 2524 39980
rect 240 39790 2524 39824
rect 240 39634 2524 39668
rect 240 39478 2524 39512
rect 240 39322 2524 39356
rect 240 39166 2524 39200
rect 240 39010 2524 39044
rect 240 38854 2524 38888
rect 240 38698 2524 38732
rect 240 38542 2524 38576
rect 240 38386 2524 38420
rect 240 38230 2524 38264
rect 240 38074 2524 38108
rect 240 37918 2524 37952
rect 240 37762 2524 37796
rect 240 37606 2524 37640
rect 240 37450 2524 37484
rect 240 37294 2524 37328
rect 240 37138 2524 37172
rect 240 36982 2524 37016
rect 240 36826 2524 36860
rect 240 36670 2524 36704
rect 240 36514 2524 36548
rect 240 36358 2524 36392
rect 240 36202 2524 36236
rect 240 36046 2524 36080
rect 240 35890 2524 35924
rect 240 35734 2524 35768
rect 240 35578 2524 35612
rect 240 35422 2524 35456
rect 240 35266 2524 35300
rect 240 35110 2524 35144
rect 240 34954 2524 34988
rect 240 34798 2524 34832
rect 240 34642 2524 34676
rect 240 34486 2524 34520
rect 240 34330 2524 34364
rect 240 34174 2524 34208
rect 240 34018 2524 34052
rect 240 33862 2524 33896
rect 240 33706 2524 33740
rect 240 33550 2524 33584
rect 240 33394 2524 33428
rect 240 33238 2524 33272
rect 240 33082 2524 33116
rect 240 32926 2524 32960
rect 240 32770 2524 32804
rect 240 32614 2524 32648
rect 240 32458 2524 32492
rect 240 32302 2524 32336
rect 240 32146 2524 32180
rect 240 31990 2524 32024
rect 240 31834 2524 31868
rect 240 31678 2524 31712
rect 240 31522 2524 31556
rect 240 31366 2524 31400
rect 240 31210 2524 31244
rect 240 31054 2524 31088
rect 240 30898 2524 30932
rect 240 30742 2524 30776
rect 240 30586 2524 30620
rect 240 30430 2524 30464
rect 240 30274 2524 30308
rect 240 30118 2524 30152
rect 240 29962 2524 29996
rect 240 29806 2524 29840
rect 240 29650 2524 29684
rect 240 29494 2524 29528
rect 240 29338 2524 29372
rect 240 29182 2524 29216
rect 240 29026 2524 29060
rect 240 28870 2524 28904
rect 240 28714 2524 28748
rect 240 28558 2524 28592
rect 240 28402 2524 28436
rect 240 28246 2524 28280
rect 240 28090 2524 28124
rect 240 27934 2524 27968
rect 240 27778 2524 27812
rect 240 27622 2524 27656
rect 240 27466 2524 27500
rect 240 27310 2524 27344
rect 240 27154 2524 27188
rect 240 26998 2524 27032
rect 240 26842 2524 26876
rect 240 26686 2524 26720
rect 240 26530 2524 26564
rect 240 26374 2524 26408
rect 240 26218 2524 26252
rect 240 26062 2524 26096
rect 240 25906 2524 25940
rect 240 25750 2524 25784
rect 240 25594 2524 25628
rect 240 25438 2524 25472
rect 240 25282 2524 25316
rect 240 25126 2524 25160
rect 240 24970 2524 25004
rect 240 24814 2524 24848
rect 240 24658 2524 24692
rect 240 24502 2524 24536
rect 240 24346 2524 24380
rect 240 24190 2524 24224
rect 240 24034 2524 24068
rect 240 23878 2524 23912
rect 240 23722 2524 23756
rect 240 23566 2524 23600
rect 240 23410 2524 23444
rect 240 23254 2524 23288
rect 240 23098 2524 23132
rect 240 22942 2524 22976
rect 240 22786 2524 22820
rect 240 22630 2524 22664
rect 240 22474 2524 22508
rect 240 22318 2524 22352
rect 240 22162 2524 22196
rect 240 22006 2524 22040
rect 240 21850 2524 21884
rect 240 21694 2524 21728
rect 240 21538 2524 21572
rect 240 21382 2524 21416
rect 240 21226 2524 21260
rect 240 21070 2524 21104
rect 240 20914 2524 20948
rect 240 20758 2524 20792
rect 240 20602 2524 20636
rect 240 20446 2524 20480
rect 240 20290 2524 20324
rect 240 20134 2524 20168
rect 240 19978 2524 20012
rect 240 19822 2524 19856
rect 240 19666 2524 19700
rect 240 19510 2524 19544
rect 240 19354 2524 19388
rect 240 19198 2524 19232
rect 240 19042 2524 19076
rect 240 18886 2524 18920
rect 240 18730 2524 18764
rect 240 18574 2524 18608
rect 240 18418 2524 18452
rect 240 18262 2524 18296
rect 240 18106 2524 18140
rect 240 17950 2524 17984
rect 240 17794 2524 17828
rect 240 17638 2524 17672
rect 240 17482 2524 17516
rect 240 17326 2524 17360
rect 240 17170 2524 17204
rect 240 17014 2524 17048
rect 240 16858 2524 16892
rect 240 16702 2524 16736
rect 240 16546 2524 16580
rect 240 16390 2524 16424
rect 240 16234 2524 16268
rect 240 16078 2524 16112
rect 240 15922 2524 15956
rect 240 15766 2524 15800
rect 240 15610 2524 15644
rect 240 15454 2524 15488
rect 240 15298 2524 15332
rect 240 15142 2524 15176
rect 240 14986 2524 15020
rect 240 14830 2524 14864
rect 240 14674 2524 14708
rect 240 14518 2524 14552
rect 240 14362 2524 14396
rect 240 14206 2524 14240
rect 240 14050 2524 14084
rect 240 13894 2524 13928
rect 240 13738 2524 13772
rect 240 13582 2524 13616
rect 240 13426 2524 13460
rect 240 13270 2524 13304
rect 240 13114 2524 13148
rect 240 12958 2524 12992
rect 240 12802 2524 12836
rect 240 12646 2524 12680
rect 240 12490 2524 12524
rect 240 12334 2524 12368
rect 240 12178 2524 12212
rect 240 12022 2524 12056
rect 240 11866 2524 11900
rect 240 11710 2524 11744
rect 240 11554 2524 11588
rect 240 11398 2524 11432
rect 240 11242 2524 11276
rect 240 11086 2524 11120
rect 240 10930 2524 10964
rect 240 10774 2524 10808
rect 240 10618 2524 10652
rect 240 10462 2524 10496
rect 240 10306 2524 10340
rect 240 10150 2524 10184
rect 240 9994 2524 10028
rect 240 9838 2524 9872
rect 240 9682 2524 9716
rect 240 9526 2524 9560
rect 240 9370 2524 9404
rect 240 9214 2524 9248
rect 240 9058 2524 9092
rect 240 8902 2524 8936
rect 240 8746 2524 8780
rect 240 8590 2524 8624
rect 240 8434 2524 8468
rect 240 8278 2524 8312
rect 240 8122 2524 8156
rect 240 7966 2524 8000
rect 240 7810 2524 7844
rect 240 7654 2524 7688
rect 240 7498 2524 7532
rect 240 7342 2524 7376
rect 240 7186 2524 7220
rect 240 7030 2524 7064
rect 240 6874 2524 6908
rect 240 6718 2524 6752
rect 240 6562 2524 6596
rect 240 6406 2524 6440
rect 240 6250 2524 6284
rect 240 6094 2524 6128
rect 240 5938 2524 5972
rect 240 5782 2524 5816
rect 240 5626 2524 5660
rect 240 5470 2524 5504
rect 240 5314 2524 5348
rect 240 5158 2524 5192
rect 240 5002 2524 5036
rect 240 4846 2524 4880
rect 240 4690 2524 4724
rect 240 4534 2524 4568
rect 240 4378 2524 4412
rect 240 4222 2524 4256
rect 240 4066 2524 4100
rect 240 3910 2524 3944
rect 240 3754 2524 3788
rect 240 3598 2524 3632
rect 240 3442 2524 3476
rect 240 3286 2524 3320
rect 240 3130 2524 3164
rect 240 2974 2524 3008
rect 240 2818 2524 2852
rect 240 2662 2524 2696
rect 240 2506 2524 2540
rect 240 2350 2524 2384
rect 240 2194 2524 2228
rect 240 2038 2524 2072
rect 240 1882 2524 1916
rect 240 1726 2524 1760
rect 240 1570 2524 1604
rect 240 1414 2524 1448
rect 240 1258 2524 1292
rect 240 1102 2524 1136
rect 240 946 2524 980
rect 240 790 2524 824
rect 240 634 2524 668
rect 240 478 2524 512
rect 240 322 2524 356
rect 150 239 184 243
rect 240 166 2524 200
rect 2586 130 2620 42980
rect 130 66 2556 100
<< metal1 >>
rect 60 43044 2626 43050
rect 60 43010 130 43044
rect 2556 43010 2626 43044
rect 60 43004 2626 43010
rect 60 42980 106 43004
rect 60 130 66 42980
rect 100 130 106 42980
rect 2580 42980 2626 43004
rect 262 42950 268 42953
rect 228 42944 268 42950
rect 1336 42950 1342 42953
rect 1336 42944 2536 42950
rect 228 42910 240 42944
rect 2524 42910 2536 42944
rect 228 42904 268 42910
rect 262 42901 268 42904
rect 1336 42904 2536 42910
rect 1336 42901 1342 42904
rect 140 42877 194 42883
rect 1422 42794 1428 42797
rect 228 42788 1428 42794
rect 2496 42794 2502 42797
rect 2496 42788 2536 42794
rect 228 42754 240 42788
rect 2524 42754 2536 42788
rect 228 42748 1428 42754
rect 1422 42745 1428 42748
rect 2496 42748 2536 42754
rect 2496 42745 2502 42748
rect 262 42638 268 42641
rect 228 42632 268 42638
rect 1336 42638 1342 42641
rect 1336 42632 2536 42638
rect 228 42598 240 42632
rect 2524 42598 2536 42632
rect 228 42592 268 42598
rect 262 42589 268 42592
rect 1336 42592 2536 42598
rect 1336 42589 1342 42592
rect 1422 42482 1428 42485
rect 228 42476 1428 42482
rect 2496 42482 2502 42485
rect 2496 42476 2536 42482
rect 228 42442 240 42476
rect 2524 42442 2536 42476
rect 228 42436 1428 42442
rect 1422 42433 1428 42436
rect 2496 42436 2536 42442
rect 2496 42433 2502 42436
rect 262 42326 268 42329
rect 228 42320 268 42326
rect 1336 42326 1342 42329
rect 1336 42320 2536 42326
rect 228 42286 240 42320
rect 2524 42286 2536 42320
rect 228 42280 268 42286
rect 262 42277 268 42280
rect 1336 42280 2536 42286
rect 1336 42277 1342 42280
rect 1422 42170 1428 42173
rect 228 42164 1428 42170
rect 2496 42170 2502 42173
rect 2496 42164 2536 42170
rect 228 42130 240 42164
rect 2524 42130 2536 42164
rect 228 42124 1428 42130
rect 1422 42121 1428 42124
rect 2496 42124 2536 42130
rect 2496 42121 2502 42124
rect 262 42014 268 42017
rect 228 42008 268 42014
rect 1336 42014 1342 42017
rect 1336 42008 2536 42014
rect 228 41974 240 42008
rect 2524 41974 2536 42008
rect 228 41968 268 41974
rect 262 41965 268 41968
rect 1336 41968 2536 41974
rect 1336 41965 1342 41968
rect 1422 41858 1428 41861
rect 228 41852 1428 41858
rect 2496 41858 2502 41861
rect 2496 41852 2536 41858
rect 228 41818 240 41852
rect 2524 41818 2536 41852
rect 228 41812 1428 41818
rect 1422 41809 1428 41812
rect 2496 41812 2536 41818
rect 2496 41809 2502 41812
rect 262 41702 268 41705
rect 228 41696 268 41702
rect 1336 41702 1342 41705
rect 1336 41696 2536 41702
rect 228 41662 240 41696
rect 2524 41662 2536 41696
rect 228 41656 268 41662
rect 262 41653 268 41656
rect 1336 41656 2536 41662
rect 1336 41653 1342 41656
rect 1422 41546 1428 41549
rect 228 41540 1428 41546
rect 2496 41546 2502 41549
rect 2496 41540 2536 41546
rect 228 41506 240 41540
rect 2524 41506 2536 41540
rect 228 41500 1428 41506
rect 1422 41497 1428 41500
rect 2496 41500 2536 41506
rect 2496 41497 2502 41500
rect 262 41390 268 41393
rect 228 41384 268 41390
rect 1336 41390 1342 41393
rect 1336 41384 2536 41390
rect 228 41350 240 41384
rect 2524 41350 2536 41384
rect 228 41344 268 41350
rect 262 41341 268 41344
rect 1336 41344 2536 41350
rect 1336 41341 1342 41344
rect 1422 41234 1428 41237
rect 228 41228 1428 41234
rect 2496 41234 2502 41237
rect 2496 41228 2536 41234
rect 228 41194 240 41228
rect 2524 41194 2536 41228
rect 228 41188 1428 41194
rect 1422 41185 1428 41188
rect 2496 41188 2536 41194
rect 2496 41185 2502 41188
rect 262 41078 268 41081
rect 228 41072 268 41078
rect 1336 41078 1342 41081
rect 1336 41072 2536 41078
rect 228 41038 240 41072
rect 2524 41038 2536 41072
rect 228 41032 268 41038
rect 262 41029 268 41032
rect 1336 41032 2536 41038
rect 1336 41029 1342 41032
rect 1422 40922 1428 40925
rect 228 40916 1428 40922
rect 2496 40922 2502 40925
rect 2496 40916 2536 40922
rect 228 40882 240 40916
rect 2524 40882 2536 40916
rect 228 40876 1428 40882
rect 1422 40873 1428 40876
rect 2496 40876 2536 40882
rect 2496 40873 2502 40876
rect 262 40766 268 40769
rect 228 40760 268 40766
rect 1336 40766 1342 40769
rect 1336 40760 2536 40766
rect 228 40726 240 40760
rect 2524 40726 2536 40760
rect 228 40720 268 40726
rect 262 40717 268 40720
rect 1336 40720 2536 40726
rect 1336 40717 1342 40720
rect 1422 40610 1428 40613
rect 228 40604 1428 40610
rect 2496 40610 2502 40613
rect 2496 40604 2536 40610
rect 228 40570 240 40604
rect 2524 40570 2536 40604
rect 228 40564 1428 40570
rect 1422 40561 1428 40564
rect 2496 40564 2536 40570
rect 2496 40561 2502 40564
rect 262 40454 268 40457
rect 228 40448 268 40454
rect 1336 40454 1342 40457
rect 1336 40448 2536 40454
rect 228 40414 240 40448
rect 2524 40414 2536 40448
rect 228 40408 268 40414
rect 262 40405 268 40408
rect 1336 40408 2536 40414
rect 1336 40405 1342 40408
rect 1422 40298 1428 40301
rect 228 40292 1428 40298
rect 2496 40298 2502 40301
rect 2496 40292 2536 40298
rect 228 40258 240 40292
rect 2524 40258 2536 40292
rect 228 40252 1428 40258
rect 1422 40249 1428 40252
rect 2496 40252 2536 40258
rect 2496 40249 2502 40252
rect 262 40142 268 40145
rect 228 40136 268 40142
rect 1336 40142 1342 40145
rect 1336 40136 2536 40142
rect 228 40102 240 40136
rect 2524 40102 2536 40136
rect 228 40096 268 40102
rect 262 40093 268 40096
rect 1336 40096 2536 40102
rect 1336 40093 1342 40096
rect 1422 39986 1428 39989
rect 228 39980 1428 39986
rect 2496 39986 2502 39989
rect 2496 39980 2536 39986
rect 228 39946 240 39980
rect 2524 39946 2536 39980
rect 228 39940 1428 39946
rect 1422 39937 1428 39940
rect 2496 39940 2536 39946
rect 2496 39937 2502 39940
rect 262 39830 268 39833
rect 228 39824 268 39830
rect 1336 39830 1342 39833
rect 1336 39824 2536 39830
rect 228 39790 240 39824
rect 2524 39790 2536 39824
rect 228 39784 268 39790
rect 262 39781 268 39784
rect 1336 39784 2536 39790
rect 1336 39781 1342 39784
rect 1422 39674 1428 39677
rect 228 39668 1428 39674
rect 2496 39674 2502 39677
rect 2496 39668 2536 39674
rect 228 39634 240 39668
rect 2524 39634 2536 39668
rect 228 39628 1428 39634
rect 1422 39625 1428 39628
rect 2496 39628 2536 39634
rect 2496 39625 2502 39628
rect 262 39518 268 39521
rect 228 39512 268 39518
rect 1336 39518 1342 39521
rect 1336 39512 2536 39518
rect 228 39478 240 39512
rect 2524 39478 2536 39512
rect 228 39472 268 39478
rect 262 39469 268 39472
rect 1336 39472 2536 39478
rect 1336 39469 1342 39472
rect 1422 39362 1428 39365
rect 228 39356 1428 39362
rect 2496 39362 2502 39365
rect 2496 39356 2536 39362
rect 228 39322 240 39356
rect 2524 39322 2536 39356
rect 228 39316 1428 39322
rect 1422 39313 1428 39316
rect 2496 39316 2536 39322
rect 2496 39313 2502 39316
rect 262 39206 268 39209
rect 228 39200 268 39206
rect 1336 39206 1342 39209
rect 1336 39200 2536 39206
rect 228 39166 240 39200
rect 2524 39166 2536 39200
rect 228 39160 268 39166
rect 262 39157 268 39160
rect 1336 39160 2536 39166
rect 1336 39157 1342 39160
rect 1422 39050 1428 39053
rect 228 39044 1428 39050
rect 2496 39050 2502 39053
rect 2496 39044 2536 39050
rect 228 39010 240 39044
rect 2524 39010 2536 39044
rect 228 39004 1428 39010
rect 1422 39001 1428 39004
rect 2496 39004 2536 39010
rect 2496 39001 2502 39004
rect 262 38894 268 38897
rect 228 38888 268 38894
rect 1336 38894 1342 38897
rect 1336 38888 2536 38894
rect 228 38854 240 38888
rect 2524 38854 2536 38888
rect 228 38848 268 38854
rect 262 38845 268 38848
rect 1336 38848 2536 38854
rect 1336 38845 1342 38848
rect 1422 38738 1428 38741
rect 228 38732 1428 38738
rect 2496 38738 2502 38741
rect 2496 38732 2536 38738
rect 228 38698 240 38732
rect 2524 38698 2536 38732
rect 228 38692 1428 38698
rect 1422 38689 1428 38692
rect 2496 38692 2536 38698
rect 2496 38689 2502 38692
rect 262 38582 268 38585
rect 228 38576 268 38582
rect 1336 38582 1342 38585
rect 1336 38576 2536 38582
rect 228 38542 240 38576
rect 2524 38542 2536 38576
rect 228 38536 268 38542
rect 262 38533 268 38536
rect 1336 38536 2536 38542
rect 1336 38533 1342 38536
rect 1422 38426 1428 38429
rect 228 38420 1428 38426
rect 2496 38426 2502 38429
rect 2496 38420 2536 38426
rect 228 38386 240 38420
rect 2524 38386 2536 38420
rect 228 38380 1428 38386
rect 1422 38377 1428 38380
rect 2496 38380 2536 38386
rect 2496 38377 2502 38380
rect 262 38270 268 38273
rect 228 38264 268 38270
rect 1336 38270 1342 38273
rect 1336 38264 2536 38270
rect 228 38230 240 38264
rect 2524 38230 2536 38264
rect 228 38224 268 38230
rect 262 38221 268 38224
rect 1336 38224 2536 38230
rect 1336 38221 1342 38224
rect 1422 38114 1428 38117
rect 228 38108 1428 38114
rect 2496 38114 2502 38117
rect 2496 38108 2536 38114
rect 228 38074 240 38108
rect 2524 38074 2536 38108
rect 228 38068 1428 38074
rect 1422 38065 1428 38068
rect 2496 38068 2536 38074
rect 2496 38065 2502 38068
rect 262 37958 268 37961
rect 228 37952 268 37958
rect 1336 37958 1342 37961
rect 1336 37952 2536 37958
rect 228 37918 240 37952
rect 2524 37918 2536 37952
rect 228 37912 268 37918
rect 262 37909 268 37912
rect 1336 37912 2536 37918
rect 1336 37909 1342 37912
rect 1422 37802 1428 37805
rect 228 37796 1428 37802
rect 2496 37802 2502 37805
rect 2496 37796 2536 37802
rect 228 37762 240 37796
rect 2524 37762 2536 37796
rect 228 37756 1428 37762
rect 1422 37753 1428 37756
rect 2496 37756 2536 37762
rect 2496 37753 2502 37756
rect 262 37646 268 37649
rect 228 37640 268 37646
rect 1336 37646 1342 37649
rect 1336 37640 2536 37646
rect 228 37606 240 37640
rect 2524 37606 2536 37640
rect 228 37600 268 37606
rect 262 37597 268 37600
rect 1336 37600 2536 37606
rect 1336 37597 1342 37600
rect 1422 37490 1428 37493
rect 228 37484 1428 37490
rect 2496 37490 2502 37493
rect 2496 37484 2536 37490
rect 228 37450 240 37484
rect 2524 37450 2536 37484
rect 228 37444 1428 37450
rect 1422 37441 1428 37444
rect 2496 37444 2536 37450
rect 2496 37441 2502 37444
rect 262 37334 268 37337
rect 228 37328 268 37334
rect 1336 37334 1342 37337
rect 1336 37328 2536 37334
rect 228 37294 240 37328
rect 2524 37294 2536 37328
rect 228 37288 268 37294
rect 262 37285 268 37288
rect 1336 37288 2536 37294
rect 1336 37285 1342 37288
rect 1422 37178 1428 37181
rect 228 37172 1428 37178
rect 2496 37178 2502 37181
rect 2496 37172 2536 37178
rect 228 37138 240 37172
rect 2524 37138 2536 37172
rect 228 37132 1428 37138
rect 1422 37129 1428 37132
rect 2496 37132 2536 37138
rect 2496 37129 2502 37132
rect 262 37022 268 37025
rect 228 37016 268 37022
rect 1336 37022 1342 37025
rect 1336 37016 2536 37022
rect 228 36982 240 37016
rect 2524 36982 2536 37016
rect 228 36976 268 36982
rect 262 36973 268 36976
rect 1336 36976 2536 36982
rect 1336 36973 1342 36976
rect 1422 36866 1428 36869
rect 228 36860 1428 36866
rect 2496 36866 2502 36869
rect 2496 36860 2536 36866
rect 228 36826 240 36860
rect 2524 36826 2536 36860
rect 228 36820 1428 36826
rect 1422 36817 1428 36820
rect 2496 36820 2536 36826
rect 2496 36817 2502 36820
rect 262 36710 268 36713
rect 228 36704 268 36710
rect 1336 36710 1342 36713
rect 1336 36704 2536 36710
rect 228 36670 240 36704
rect 2524 36670 2536 36704
rect 228 36664 268 36670
rect 262 36661 268 36664
rect 1336 36664 2536 36670
rect 1336 36661 1342 36664
rect 1422 36554 1428 36557
rect 228 36548 1428 36554
rect 2496 36554 2502 36557
rect 2496 36548 2536 36554
rect 228 36514 240 36548
rect 2524 36514 2536 36548
rect 228 36508 1428 36514
rect 1422 36505 1428 36508
rect 2496 36508 2536 36514
rect 2496 36505 2502 36508
rect 262 36398 268 36401
rect 228 36392 268 36398
rect 1336 36398 1342 36401
rect 1336 36392 2536 36398
rect 228 36358 240 36392
rect 2524 36358 2536 36392
rect 228 36352 268 36358
rect 262 36349 268 36352
rect 1336 36352 2536 36358
rect 1336 36349 1342 36352
rect 1422 36242 1428 36245
rect 228 36236 1428 36242
rect 2496 36242 2502 36245
rect 2496 36236 2536 36242
rect 228 36202 240 36236
rect 2524 36202 2536 36236
rect 228 36196 1428 36202
rect 1422 36193 1428 36196
rect 2496 36196 2536 36202
rect 2496 36193 2502 36196
rect 262 36086 268 36089
rect 228 36080 268 36086
rect 1336 36086 1342 36089
rect 1336 36080 2536 36086
rect 228 36046 240 36080
rect 2524 36046 2536 36080
rect 228 36040 268 36046
rect 262 36037 268 36040
rect 1336 36040 2536 36046
rect 1336 36037 1342 36040
rect 1422 35930 1428 35933
rect 228 35924 1428 35930
rect 2496 35930 2502 35933
rect 2496 35924 2536 35930
rect 228 35890 240 35924
rect 2524 35890 2536 35924
rect 228 35884 1428 35890
rect 1422 35881 1428 35884
rect 2496 35884 2536 35890
rect 2496 35881 2502 35884
rect 262 35774 268 35777
rect 228 35768 268 35774
rect 1336 35774 1342 35777
rect 1336 35768 2536 35774
rect 228 35734 240 35768
rect 2524 35734 2536 35768
rect 228 35728 268 35734
rect 262 35725 268 35728
rect 1336 35728 2536 35734
rect 1336 35725 1342 35728
rect 1422 35618 1428 35621
rect 228 35612 1428 35618
rect 2496 35618 2502 35621
rect 2496 35612 2536 35618
rect 228 35578 240 35612
rect 2524 35578 2536 35612
rect 228 35572 1428 35578
rect 1422 35569 1428 35572
rect 2496 35572 2536 35578
rect 2496 35569 2502 35572
rect 262 35462 268 35465
rect 228 35456 268 35462
rect 1336 35462 1342 35465
rect 1336 35456 2536 35462
rect 228 35422 240 35456
rect 2524 35422 2536 35456
rect 228 35416 268 35422
rect 262 35413 268 35416
rect 1336 35416 2536 35422
rect 1336 35413 1342 35416
rect 1422 35306 1428 35309
rect 228 35300 1428 35306
rect 2496 35306 2502 35309
rect 2496 35300 2536 35306
rect 228 35266 240 35300
rect 2524 35266 2536 35300
rect 228 35260 1428 35266
rect 1422 35257 1428 35260
rect 2496 35260 2536 35266
rect 2496 35257 2502 35260
rect 262 35150 268 35153
rect 228 35144 268 35150
rect 1336 35150 1342 35153
rect 1336 35144 2536 35150
rect 228 35110 240 35144
rect 2524 35110 2536 35144
rect 228 35104 268 35110
rect 262 35101 268 35104
rect 1336 35104 2536 35110
rect 1336 35101 1342 35104
rect 1422 34994 1428 34997
rect 228 34988 1428 34994
rect 2496 34994 2502 34997
rect 2496 34988 2536 34994
rect 228 34954 240 34988
rect 2524 34954 2536 34988
rect 228 34948 1428 34954
rect 1422 34945 1428 34948
rect 2496 34948 2536 34954
rect 2496 34945 2502 34948
rect 262 34838 268 34841
rect 228 34832 268 34838
rect 1336 34838 1342 34841
rect 1336 34832 2536 34838
rect 228 34798 240 34832
rect 2524 34798 2536 34832
rect 228 34792 268 34798
rect 262 34789 268 34792
rect 1336 34792 2536 34798
rect 1336 34789 1342 34792
rect 1422 34682 1428 34685
rect 228 34676 1428 34682
rect 2496 34682 2502 34685
rect 2496 34676 2536 34682
rect 228 34642 240 34676
rect 2524 34642 2536 34676
rect 228 34636 1428 34642
rect 1422 34633 1428 34636
rect 2496 34636 2536 34642
rect 2496 34633 2502 34636
rect 262 34526 268 34529
rect 228 34520 268 34526
rect 1336 34526 1342 34529
rect 1336 34520 2536 34526
rect 228 34486 240 34520
rect 2524 34486 2536 34520
rect 228 34480 268 34486
rect 262 34477 268 34480
rect 1336 34480 2536 34486
rect 1336 34477 1342 34480
rect 1422 34370 1428 34373
rect 228 34364 1428 34370
rect 2496 34370 2502 34373
rect 2496 34364 2536 34370
rect 228 34330 240 34364
rect 2524 34330 2536 34364
rect 228 34324 1428 34330
rect 1422 34321 1428 34324
rect 2496 34324 2536 34330
rect 2496 34321 2502 34324
rect 262 34214 268 34217
rect 228 34208 268 34214
rect 1336 34214 1342 34217
rect 1336 34208 2536 34214
rect 228 34174 240 34208
rect 2524 34174 2536 34208
rect 228 34168 268 34174
rect 262 34165 268 34168
rect 1336 34168 2536 34174
rect 1336 34165 1342 34168
rect 1422 34058 1428 34061
rect 228 34052 1428 34058
rect 2496 34058 2502 34061
rect 2496 34052 2536 34058
rect 228 34018 240 34052
rect 2524 34018 2536 34052
rect 228 34012 1428 34018
rect 1422 34009 1428 34012
rect 2496 34012 2536 34018
rect 2496 34009 2502 34012
rect 262 33902 268 33905
rect 228 33896 268 33902
rect 1336 33902 1342 33905
rect 1336 33896 2536 33902
rect 228 33862 240 33896
rect 2524 33862 2536 33896
rect 228 33856 268 33862
rect 262 33853 268 33856
rect 1336 33856 2536 33862
rect 1336 33853 1342 33856
rect 1422 33746 1428 33749
rect 228 33740 1428 33746
rect 2496 33746 2502 33749
rect 2496 33740 2536 33746
rect 228 33706 240 33740
rect 2524 33706 2536 33740
rect 228 33700 1428 33706
rect 1422 33697 1428 33700
rect 2496 33700 2536 33706
rect 2496 33697 2502 33700
rect 262 33590 268 33593
rect 228 33584 268 33590
rect 1336 33590 1342 33593
rect 1336 33584 2536 33590
rect 228 33550 240 33584
rect 2524 33550 2536 33584
rect 228 33544 268 33550
rect 262 33541 268 33544
rect 1336 33544 2536 33550
rect 1336 33541 1342 33544
rect 1422 33434 1428 33437
rect 228 33428 1428 33434
rect 2496 33434 2502 33437
rect 2496 33428 2536 33434
rect 228 33394 240 33428
rect 2524 33394 2536 33428
rect 228 33388 1428 33394
rect 1422 33385 1428 33388
rect 2496 33388 2536 33394
rect 2496 33385 2502 33388
rect 262 33278 268 33281
rect 228 33272 268 33278
rect 1336 33278 1342 33281
rect 1336 33272 2536 33278
rect 228 33238 240 33272
rect 2524 33238 2536 33272
rect 228 33232 268 33238
rect 262 33229 268 33232
rect 1336 33232 2536 33238
rect 1336 33229 1342 33232
rect 1422 33122 1428 33125
rect 228 33116 1428 33122
rect 2496 33122 2502 33125
rect 2496 33116 2536 33122
rect 228 33082 240 33116
rect 2524 33082 2536 33116
rect 228 33076 1428 33082
rect 1422 33073 1428 33076
rect 2496 33076 2536 33082
rect 2496 33073 2502 33076
rect 262 32966 268 32969
rect 228 32960 268 32966
rect 1336 32966 1342 32969
rect 1336 32960 2536 32966
rect 228 32926 240 32960
rect 2524 32926 2536 32960
rect 228 32920 268 32926
rect 262 32917 268 32920
rect 1336 32920 2536 32926
rect 1336 32917 1342 32920
rect 1422 32810 1428 32813
rect 228 32804 1428 32810
rect 2496 32810 2502 32813
rect 2496 32804 2536 32810
rect 228 32770 240 32804
rect 2524 32770 2536 32804
rect 228 32764 1428 32770
rect 1422 32761 1428 32764
rect 2496 32764 2536 32770
rect 2496 32761 2502 32764
rect 262 32654 268 32657
rect 228 32648 268 32654
rect 1336 32654 1342 32657
rect 1336 32648 2536 32654
rect 228 32614 240 32648
rect 2524 32614 2536 32648
rect 228 32608 268 32614
rect 262 32605 268 32608
rect 1336 32608 2536 32614
rect 1336 32605 1342 32608
rect 1422 32498 1428 32501
rect 228 32492 1428 32498
rect 2496 32498 2502 32501
rect 2496 32492 2536 32498
rect 228 32458 240 32492
rect 2524 32458 2536 32492
rect 228 32452 1428 32458
rect 1422 32449 1428 32452
rect 2496 32452 2536 32458
rect 2496 32449 2502 32452
rect 262 32342 268 32345
rect 228 32336 268 32342
rect 1336 32342 1342 32345
rect 1336 32336 2536 32342
rect 228 32302 240 32336
rect 2524 32302 2536 32336
rect 228 32296 268 32302
rect 262 32293 268 32296
rect 1336 32296 2536 32302
rect 1336 32293 1342 32296
rect 1422 32186 1428 32189
rect 228 32180 1428 32186
rect 2496 32186 2502 32189
rect 2496 32180 2536 32186
rect 228 32146 240 32180
rect 2524 32146 2536 32180
rect 228 32140 1428 32146
rect 1422 32137 1428 32140
rect 2496 32140 2536 32146
rect 2496 32137 2502 32140
rect 262 32030 268 32033
rect 228 32024 268 32030
rect 1336 32030 1342 32033
rect 1336 32024 2536 32030
rect 228 31990 240 32024
rect 2524 31990 2536 32024
rect 228 31984 268 31990
rect 262 31981 268 31984
rect 1336 31984 2536 31990
rect 1336 31981 1342 31984
rect 1422 31874 1428 31877
rect 228 31868 1428 31874
rect 2496 31874 2502 31877
rect 2496 31868 2536 31874
rect 228 31834 240 31868
rect 2524 31834 2536 31868
rect 228 31828 1428 31834
rect 1422 31825 1428 31828
rect 2496 31828 2536 31834
rect 2496 31825 2502 31828
rect 262 31718 268 31721
rect 228 31712 268 31718
rect 1336 31718 1342 31721
rect 1336 31712 2536 31718
rect 228 31678 240 31712
rect 2524 31678 2536 31712
rect 228 31672 268 31678
rect 262 31669 268 31672
rect 1336 31672 2536 31678
rect 1336 31669 1342 31672
rect 1422 31562 1428 31565
rect 228 31556 1428 31562
rect 2496 31562 2502 31565
rect 2496 31556 2536 31562
rect 228 31522 240 31556
rect 2524 31522 2536 31556
rect 228 31516 1428 31522
rect 1422 31513 1428 31516
rect 2496 31516 2536 31522
rect 2496 31513 2502 31516
rect 262 31406 268 31409
rect 228 31400 268 31406
rect 1336 31406 1342 31409
rect 1336 31400 2536 31406
rect 228 31366 240 31400
rect 2524 31366 2536 31400
rect 228 31360 268 31366
rect 262 31357 268 31360
rect 1336 31360 2536 31366
rect 1336 31357 1342 31360
rect 1422 31250 1428 31253
rect 228 31244 1428 31250
rect 2496 31250 2502 31253
rect 2496 31244 2536 31250
rect 228 31210 240 31244
rect 2524 31210 2536 31244
rect 228 31204 1428 31210
rect 1422 31201 1428 31204
rect 2496 31204 2536 31210
rect 2496 31201 2502 31204
rect 262 31094 268 31097
rect 228 31088 268 31094
rect 1336 31094 1342 31097
rect 1336 31088 2536 31094
rect 228 31054 240 31088
rect 2524 31054 2536 31088
rect 228 31048 268 31054
rect 262 31045 268 31048
rect 1336 31048 2536 31054
rect 1336 31045 1342 31048
rect 1422 30938 1428 30941
rect 228 30932 1428 30938
rect 2496 30938 2502 30941
rect 2496 30932 2536 30938
rect 228 30898 240 30932
rect 2524 30898 2536 30932
rect 228 30892 1428 30898
rect 1422 30889 1428 30892
rect 2496 30892 2536 30898
rect 2496 30889 2502 30892
rect 262 30782 268 30785
rect 228 30776 268 30782
rect 1336 30782 1342 30785
rect 1336 30776 2536 30782
rect 228 30742 240 30776
rect 2524 30742 2536 30776
rect 228 30736 268 30742
rect 262 30733 268 30736
rect 1336 30736 2536 30742
rect 1336 30733 1342 30736
rect 1422 30626 1428 30629
rect 228 30620 1428 30626
rect 2496 30626 2502 30629
rect 2496 30620 2536 30626
rect 228 30586 240 30620
rect 2524 30586 2536 30620
rect 228 30580 1428 30586
rect 1422 30577 1428 30580
rect 2496 30580 2536 30586
rect 2496 30577 2502 30580
rect 262 30470 268 30473
rect 228 30464 268 30470
rect 1336 30470 1342 30473
rect 1336 30464 2536 30470
rect 228 30430 240 30464
rect 2524 30430 2536 30464
rect 228 30424 268 30430
rect 262 30421 268 30424
rect 1336 30424 2536 30430
rect 1336 30421 1342 30424
rect 1422 30314 1428 30317
rect 228 30308 1428 30314
rect 2496 30314 2502 30317
rect 2496 30308 2536 30314
rect 228 30274 240 30308
rect 2524 30274 2536 30308
rect 228 30268 1428 30274
rect 1422 30265 1428 30268
rect 2496 30268 2536 30274
rect 2496 30265 2502 30268
rect 262 30158 268 30161
rect 228 30152 268 30158
rect 1336 30158 1342 30161
rect 1336 30152 2536 30158
rect 228 30118 240 30152
rect 2524 30118 2536 30152
rect 228 30112 268 30118
rect 262 30109 268 30112
rect 1336 30112 2536 30118
rect 1336 30109 1342 30112
rect 1422 30002 1428 30005
rect 228 29996 1428 30002
rect 2496 30002 2502 30005
rect 2496 29996 2536 30002
rect 228 29962 240 29996
rect 2524 29962 2536 29996
rect 228 29956 1428 29962
rect 1422 29953 1428 29956
rect 2496 29956 2536 29962
rect 2496 29953 2502 29956
rect 262 29846 268 29849
rect 228 29840 268 29846
rect 1336 29846 1342 29849
rect 1336 29840 2536 29846
rect 228 29806 240 29840
rect 2524 29806 2536 29840
rect 228 29800 268 29806
rect 262 29797 268 29800
rect 1336 29800 2536 29806
rect 1336 29797 1342 29800
rect 1422 29690 1428 29693
rect 228 29684 1428 29690
rect 2496 29690 2502 29693
rect 2496 29684 2536 29690
rect 228 29650 240 29684
rect 2524 29650 2536 29684
rect 228 29644 1428 29650
rect 1422 29641 1428 29644
rect 2496 29644 2536 29650
rect 2496 29641 2502 29644
rect 262 29534 268 29537
rect 228 29528 268 29534
rect 1336 29534 1342 29537
rect 1336 29528 2536 29534
rect 228 29494 240 29528
rect 2524 29494 2536 29528
rect 228 29488 268 29494
rect 262 29485 268 29488
rect 1336 29488 2536 29494
rect 1336 29485 1342 29488
rect 1422 29378 1428 29381
rect 228 29372 1428 29378
rect 2496 29378 2502 29381
rect 2496 29372 2536 29378
rect 228 29338 240 29372
rect 2524 29338 2536 29372
rect 228 29332 1428 29338
rect 1422 29329 1428 29332
rect 2496 29332 2536 29338
rect 2496 29329 2502 29332
rect 262 29222 268 29225
rect 228 29216 268 29222
rect 1336 29222 1342 29225
rect 1336 29216 2536 29222
rect 228 29182 240 29216
rect 2524 29182 2536 29216
rect 228 29176 268 29182
rect 262 29173 268 29176
rect 1336 29176 2536 29182
rect 1336 29173 1342 29176
rect 1422 29066 1428 29069
rect 228 29060 1428 29066
rect 2496 29066 2502 29069
rect 2496 29060 2536 29066
rect 228 29026 240 29060
rect 2524 29026 2536 29060
rect 228 29020 1428 29026
rect 1422 29017 1428 29020
rect 2496 29020 2536 29026
rect 2496 29017 2502 29020
rect 262 28910 268 28913
rect 228 28904 268 28910
rect 1336 28910 1342 28913
rect 1336 28904 2536 28910
rect 228 28870 240 28904
rect 2524 28870 2536 28904
rect 228 28864 268 28870
rect 262 28861 268 28864
rect 1336 28864 2536 28870
rect 1336 28861 1342 28864
rect 1422 28754 1428 28757
rect 228 28748 1428 28754
rect 2496 28754 2502 28757
rect 2496 28748 2536 28754
rect 228 28714 240 28748
rect 2524 28714 2536 28748
rect 228 28708 1428 28714
rect 1422 28705 1428 28708
rect 2496 28708 2536 28714
rect 2496 28705 2502 28708
rect 262 28598 268 28601
rect 228 28592 268 28598
rect 1336 28598 1342 28601
rect 1336 28592 2536 28598
rect 228 28558 240 28592
rect 2524 28558 2536 28592
rect 228 28552 268 28558
rect 262 28549 268 28552
rect 1336 28552 2536 28558
rect 1336 28549 1342 28552
rect 1422 28442 1428 28445
rect 228 28436 1428 28442
rect 2496 28442 2502 28445
rect 2496 28436 2536 28442
rect 228 28402 240 28436
rect 2524 28402 2536 28436
rect 228 28396 1428 28402
rect 1422 28393 1428 28396
rect 2496 28396 2536 28402
rect 2496 28393 2502 28396
rect 262 28286 268 28289
rect 228 28280 268 28286
rect 1336 28286 1342 28289
rect 1336 28280 2536 28286
rect 228 28246 240 28280
rect 2524 28246 2536 28280
rect 228 28240 268 28246
rect 262 28237 268 28240
rect 1336 28240 2536 28246
rect 1336 28237 1342 28240
rect 1422 28130 1428 28133
rect 228 28124 1428 28130
rect 2496 28130 2502 28133
rect 2496 28124 2536 28130
rect 228 28090 240 28124
rect 2524 28090 2536 28124
rect 228 28084 1428 28090
rect 1422 28081 1428 28084
rect 2496 28084 2536 28090
rect 2496 28081 2502 28084
rect 262 27974 268 27977
rect 228 27968 268 27974
rect 1336 27974 1342 27977
rect 1336 27968 2536 27974
rect 228 27934 240 27968
rect 2524 27934 2536 27968
rect 228 27928 268 27934
rect 262 27925 268 27928
rect 1336 27928 2536 27934
rect 1336 27925 1342 27928
rect 1422 27818 1428 27821
rect 228 27812 1428 27818
rect 2496 27818 2502 27821
rect 2496 27812 2536 27818
rect 228 27778 240 27812
rect 2524 27778 2536 27812
rect 228 27772 1428 27778
rect 1422 27769 1428 27772
rect 2496 27772 2536 27778
rect 2496 27769 2502 27772
rect 262 27662 268 27665
rect 228 27656 268 27662
rect 1336 27662 1342 27665
rect 1336 27656 2536 27662
rect 228 27622 240 27656
rect 2524 27622 2536 27656
rect 228 27616 268 27622
rect 262 27613 268 27616
rect 1336 27616 2536 27622
rect 1336 27613 1342 27616
rect 1422 27506 1428 27509
rect 228 27500 1428 27506
rect 2496 27506 2502 27509
rect 2496 27500 2536 27506
rect 228 27466 240 27500
rect 2524 27466 2536 27500
rect 228 27460 1428 27466
rect 1422 27457 1428 27460
rect 2496 27460 2536 27466
rect 2496 27457 2502 27460
rect 262 27350 268 27353
rect 228 27344 268 27350
rect 1336 27350 1342 27353
rect 1336 27344 2536 27350
rect 228 27310 240 27344
rect 2524 27310 2536 27344
rect 228 27304 268 27310
rect 262 27301 268 27304
rect 1336 27304 2536 27310
rect 1336 27301 1342 27304
rect 1422 27194 1428 27197
rect 228 27188 1428 27194
rect 2496 27194 2502 27197
rect 2496 27188 2536 27194
rect 228 27154 240 27188
rect 2524 27154 2536 27188
rect 228 27148 1428 27154
rect 1422 27145 1428 27148
rect 2496 27148 2536 27154
rect 2496 27145 2502 27148
rect 262 27038 268 27041
rect 228 27032 268 27038
rect 1336 27038 1342 27041
rect 1336 27032 2536 27038
rect 228 26998 240 27032
rect 2524 26998 2536 27032
rect 228 26992 268 26998
rect 262 26989 268 26992
rect 1336 26992 2536 26998
rect 1336 26989 1342 26992
rect 1422 26882 1428 26885
rect 228 26876 1428 26882
rect 2496 26882 2502 26885
rect 2496 26876 2536 26882
rect 228 26842 240 26876
rect 2524 26842 2536 26876
rect 228 26836 1428 26842
rect 1422 26833 1428 26836
rect 2496 26836 2536 26842
rect 2496 26833 2502 26836
rect 262 26726 268 26729
rect 228 26720 268 26726
rect 1336 26726 1342 26729
rect 1336 26720 2536 26726
rect 228 26686 240 26720
rect 2524 26686 2536 26720
rect 228 26680 268 26686
rect 262 26677 268 26680
rect 1336 26680 2536 26686
rect 1336 26677 1342 26680
rect 1422 26570 1428 26573
rect 228 26564 1428 26570
rect 2496 26570 2502 26573
rect 2496 26564 2536 26570
rect 228 26530 240 26564
rect 2524 26530 2536 26564
rect 228 26524 1428 26530
rect 1422 26521 1428 26524
rect 2496 26524 2536 26530
rect 2496 26521 2502 26524
rect 262 26414 268 26417
rect 228 26408 268 26414
rect 1336 26414 1342 26417
rect 1336 26408 2536 26414
rect 228 26374 240 26408
rect 2524 26374 2536 26408
rect 228 26368 268 26374
rect 262 26365 268 26368
rect 1336 26368 2536 26374
rect 1336 26365 1342 26368
rect 1422 26258 1428 26261
rect 228 26252 1428 26258
rect 2496 26258 2502 26261
rect 2496 26252 2536 26258
rect 228 26218 240 26252
rect 2524 26218 2536 26252
rect 228 26212 1428 26218
rect 1422 26209 1428 26212
rect 2496 26212 2536 26218
rect 2496 26209 2502 26212
rect 262 26102 268 26105
rect 228 26096 268 26102
rect 1336 26102 1342 26105
rect 1336 26096 2536 26102
rect 228 26062 240 26096
rect 2524 26062 2536 26096
rect 228 26056 268 26062
rect 262 26053 268 26056
rect 1336 26056 2536 26062
rect 1336 26053 1342 26056
rect 1422 25946 1428 25949
rect 228 25940 1428 25946
rect 2496 25946 2502 25949
rect 2496 25940 2536 25946
rect 228 25906 240 25940
rect 2524 25906 2536 25940
rect 228 25900 1428 25906
rect 1422 25897 1428 25900
rect 2496 25900 2536 25906
rect 2496 25897 2502 25900
rect 262 25790 268 25793
rect 228 25784 268 25790
rect 1336 25790 1342 25793
rect 1336 25784 2536 25790
rect 228 25750 240 25784
rect 2524 25750 2536 25784
rect 228 25744 268 25750
rect 262 25741 268 25744
rect 1336 25744 2536 25750
rect 1336 25741 1342 25744
rect 1422 25634 1428 25637
rect 228 25628 1428 25634
rect 2496 25634 2502 25637
rect 2496 25628 2536 25634
rect 228 25594 240 25628
rect 2524 25594 2536 25628
rect 228 25588 1428 25594
rect 1422 25585 1428 25588
rect 2496 25588 2536 25594
rect 2496 25585 2502 25588
rect 262 25478 268 25481
rect 228 25472 268 25478
rect 1336 25478 1342 25481
rect 1336 25472 2536 25478
rect 228 25438 240 25472
rect 2524 25438 2536 25472
rect 228 25432 268 25438
rect 262 25429 268 25432
rect 1336 25432 2536 25438
rect 1336 25429 1342 25432
rect 1422 25322 1428 25325
rect 228 25316 1428 25322
rect 2496 25322 2502 25325
rect 2496 25316 2536 25322
rect 228 25282 240 25316
rect 2524 25282 2536 25316
rect 228 25276 1428 25282
rect 1422 25273 1428 25276
rect 2496 25276 2536 25282
rect 2496 25273 2502 25276
rect 262 25166 268 25169
rect 228 25160 268 25166
rect 1336 25166 1342 25169
rect 1336 25160 2536 25166
rect 228 25126 240 25160
rect 2524 25126 2536 25160
rect 228 25120 268 25126
rect 262 25117 268 25120
rect 1336 25120 2536 25126
rect 1336 25117 1342 25120
rect 1422 25010 1428 25013
rect 228 25004 1428 25010
rect 2496 25010 2502 25013
rect 2496 25004 2536 25010
rect 228 24970 240 25004
rect 2524 24970 2536 25004
rect 228 24964 1428 24970
rect 1422 24961 1428 24964
rect 2496 24964 2536 24970
rect 2496 24961 2502 24964
rect 262 24854 268 24857
rect 228 24848 268 24854
rect 1336 24854 1342 24857
rect 1336 24848 2536 24854
rect 228 24814 240 24848
rect 2524 24814 2536 24848
rect 228 24808 268 24814
rect 262 24805 268 24808
rect 1336 24808 2536 24814
rect 1336 24805 1342 24808
rect 1422 24698 1428 24701
rect 228 24692 1428 24698
rect 2496 24698 2502 24701
rect 2496 24692 2536 24698
rect 228 24658 240 24692
rect 2524 24658 2536 24692
rect 228 24652 1428 24658
rect 1422 24649 1428 24652
rect 2496 24652 2536 24658
rect 2496 24649 2502 24652
rect 262 24542 268 24545
rect 228 24536 268 24542
rect 1336 24542 1342 24545
rect 1336 24536 2536 24542
rect 228 24502 240 24536
rect 2524 24502 2536 24536
rect 228 24496 268 24502
rect 262 24493 268 24496
rect 1336 24496 2536 24502
rect 1336 24493 1342 24496
rect 1422 24386 1428 24389
rect 228 24380 1428 24386
rect 2496 24386 2502 24389
rect 2496 24380 2536 24386
rect 228 24346 240 24380
rect 2524 24346 2536 24380
rect 228 24340 1428 24346
rect 1422 24337 1428 24340
rect 2496 24340 2536 24346
rect 2496 24337 2502 24340
rect 262 24230 268 24233
rect 228 24224 268 24230
rect 1336 24230 1342 24233
rect 1336 24224 2536 24230
rect 228 24190 240 24224
rect 2524 24190 2536 24224
rect 228 24184 268 24190
rect 262 24181 268 24184
rect 1336 24184 2536 24190
rect 1336 24181 1342 24184
rect 1422 24074 1428 24077
rect 228 24068 1428 24074
rect 2496 24074 2502 24077
rect 2496 24068 2536 24074
rect 228 24034 240 24068
rect 2524 24034 2536 24068
rect 228 24028 1428 24034
rect 1422 24025 1428 24028
rect 2496 24028 2536 24034
rect 2496 24025 2502 24028
rect 262 23918 268 23921
rect 228 23912 268 23918
rect 1336 23918 1342 23921
rect 1336 23912 2536 23918
rect 228 23878 240 23912
rect 2524 23878 2536 23912
rect 228 23872 268 23878
rect 262 23869 268 23872
rect 1336 23872 2536 23878
rect 1336 23869 1342 23872
rect 1422 23762 1428 23765
rect 228 23756 1428 23762
rect 2496 23762 2502 23765
rect 2496 23756 2536 23762
rect 228 23722 240 23756
rect 2524 23722 2536 23756
rect 228 23716 1428 23722
rect 1422 23713 1428 23716
rect 2496 23716 2536 23722
rect 2496 23713 2502 23716
rect 262 23606 268 23609
rect 228 23600 268 23606
rect 1336 23606 1342 23609
rect 1336 23600 2536 23606
rect 228 23566 240 23600
rect 2524 23566 2536 23600
rect 228 23560 268 23566
rect 262 23557 268 23560
rect 1336 23560 2536 23566
rect 1336 23557 1342 23560
rect 1422 23450 1428 23453
rect 228 23444 1428 23450
rect 2496 23450 2502 23453
rect 2496 23444 2536 23450
rect 228 23410 240 23444
rect 2524 23410 2536 23444
rect 228 23404 1428 23410
rect 1422 23401 1428 23404
rect 2496 23404 2536 23410
rect 2496 23401 2502 23404
rect 262 23294 268 23297
rect 228 23288 268 23294
rect 1336 23294 1342 23297
rect 1336 23288 2536 23294
rect 228 23254 240 23288
rect 2524 23254 2536 23288
rect 228 23248 268 23254
rect 262 23245 268 23248
rect 1336 23248 2536 23254
rect 1336 23245 1342 23248
rect 1422 23138 1428 23141
rect 228 23132 1428 23138
rect 2496 23138 2502 23141
rect 2496 23132 2536 23138
rect 228 23098 240 23132
rect 2524 23098 2536 23132
rect 228 23092 1428 23098
rect 1422 23089 1428 23092
rect 2496 23092 2536 23098
rect 2496 23089 2502 23092
rect 262 22982 268 22985
rect 228 22976 268 22982
rect 1336 22982 1342 22985
rect 1336 22976 2536 22982
rect 228 22942 240 22976
rect 2524 22942 2536 22976
rect 228 22936 268 22942
rect 262 22933 268 22936
rect 1336 22936 2536 22942
rect 1336 22933 1342 22936
rect 1422 22826 1428 22829
rect 228 22820 1428 22826
rect 2496 22826 2502 22829
rect 2496 22820 2536 22826
rect 228 22786 240 22820
rect 2524 22786 2536 22820
rect 228 22780 1428 22786
rect 1422 22777 1428 22780
rect 2496 22780 2536 22786
rect 2496 22777 2502 22780
rect 262 22670 268 22673
rect 228 22664 268 22670
rect 1336 22670 1342 22673
rect 1336 22664 2536 22670
rect 228 22630 240 22664
rect 2524 22630 2536 22664
rect 228 22624 268 22630
rect 262 22621 268 22624
rect 1336 22624 2536 22630
rect 1336 22621 1342 22624
rect 1422 22514 1428 22517
rect 228 22508 1428 22514
rect 2496 22514 2502 22517
rect 2496 22508 2536 22514
rect 228 22474 240 22508
rect 2524 22474 2536 22508
rect 228 22468 1428 22474
rect 1422 22465 1428 22468
rect 2496 22468 2536 22474
rect 2496 22465 2502 22468
rect 262 22358 268 22361
rect 228 22352 268 22358
rect 1336 22358 1342 22361
rect 1336 22352 2536 22358
rect 228 22318 240 22352
rect 2524 22318 2536 22352
rect 228 22312 268 22318
rect 262 22309 268 22312
rect 1336 22312 2536 22318
rect 1336 22309 1342 22312
rect 1422 22202 1428 22205
rect 228 22196 1428 22202
rect 2496 22202 2502 22205
rect 2496 22196 2536 22202
rect 228 22162 240 22196
rect 2524 22162 2536 22196
rect 228 22156 1428 22162
rect 1422 22153 1428 22156
rect 2496 22156 2536 22162
rect 2496 22153 2502 22156
rect 262 22046 268 22049
rect 228 22040 268 22046
rect 1336 22046 1342 22049
rect 1336 22040 2536 22046
rect 228 22006 240 22040
rect 2524 22006 2536 22040
rect 228 22000 268 22006
rect 262 21997 268 22000
rect 1336 22000 2536 22006
rect 1336 21997 1342 22000
rect 1422 21890 1428 21893
rect 228 21884 1428 21890
rect 2496 21890 2502 21893
rect 2496 21884 2536 21890
rect 228 21850 240 21884
rect 2524 21850 2536 21884
rect 228 21844 1428 21850
rect 1422 21841 1428 21844
rect 2496 21844 2536 21850
rect 2496 21841 2502 21844
rect 262 21734 268 21737
rect 228 21728 268 21734
rect 1336 21734 1342 21737
rect 1336 21728 2536 21734
rect 228 21694 240 21728
rect 2524 21694 2536 21728
rect 228 21688 268 21694
rect 262 21685 268 21688
rect 1336 21688 2536 21694
rect 1336 21685 1342 21688
rect 1422 21578 1428 21581
rect 228 21572 1428 21578
rect 2496 21578 2502 21581
rect 2496 21572 2536 21578
rect 228 21538 240 21572
rect 2524 21538 2536 21572
rect 228 21532 1428 21538
rect 1422 21529 1428 21532
rect 2496 21532 2536 21538
rect 2496 21529 2502 21532
rect 262 21422 268 21425
rect 228 21416 268 21422
rect 1336 21422 1342 21425
rect 1336 21416 2536 21422
rect 228 21382 240 21416
rect 2524 21382 2536 21416
rect 228 21376 268 21382
rect 262 21373 268 21376
rect 1336 21376 2536 21382
rect 1336 21373 1342 21376
rect 1422 21266 1428 21269
rect 228 21260 1428 21266
rect 2496 21266 2502 21269
rect 2496 21260 2536 21266
rect 228 21226 240 21260
rect 2524 21226 2536 21260
rect 228 21220 1428 21226
rect 1422 21217 1428 21220
rect 2496 21220 2536 21226
rect 2496 21217 2502 21220
rect 262 21110 268 21113
rect 228 21104 268 21110
rect 1336 21110 1342 21113
rect 1336 21104 2536 21110
rect 228 21070 240 21104
rect 2524 21070 2536 21104
rect 228 21064 268 21070
rect 262 21061 268 21064
rect 1336 21064 2536 21070
rect 1336 21061 1342 21064
rect 1422 20954 1428 20957
rect 228 20948 1428 20954
rect 2496 20954 2502 20957
rect 2496 20948 2536 20954
rect 228 20914 240 20948
rect 2524 20914 2536 20948
rect 228 20908 1428 20914
rect 1422 20905 1428 20908
rect 2496 20908 2536 20914
rect 2496 20905 2502 20908
rect 262 20798 268 20801
rect 228 20792 268 20798
rect 1336 20798 1342 20801
rect 1336 20792 2536 20798
rect 228 20758 240 20792
rect 2524 20758 2536 20792
rect 228 20752 268 20758
rect 262 20749 268 20752
rect 1336 20752 2536 20758
rect 1336 20749 1342 20752
rect 1422 20642 1428 20645
rect 228 20636 1428 20642
rect 2496 20642 2502 20645
rect 2496 20636 2536 20642
rect 228 20602 240 20636
rect 2524 20602 2536 20636
rect 228 20596 1428 20602
rect 1422 20593 1428 20596
rect 2496 20596 2536 20602
rect 2496 20593 2502 20596
rect 262 20486 268 20489
rect 228 20480 268 20486
rect 1336 20486 1342 20489
rect 1336 20480 2536 20486
rect 228 20446 240 20480
rect 2524 20446 2536 20480
rect 228 20440 268 20446
rect 262 20437 268 20440
rect 1336 20440 2536 20446
rect 1336 20437 1342 20440
rect 1422 20330 1428 20333
rect 228 20324 1428 20330
rect 2496 20330 2502 20333
rect 2496 20324 2536 20330
rect 228 20290 240 20324
rect 2524 20290 2536 20324
rect 228 20284 1428 20290
rect 1422 20281 1428 20284
rect 2496 20284 2536 20290
rect 2496 20281 2502 20284
rect 262 20174 268 20177
rect 228 20168 268 20174
rect 1336 20174 1342 20177
rect 1336 20168 2536 20174
rect 228 20134 240 20168
rect 2524 20134 2536 20168
rect 228 20128 268 20134
rect 262 20125 268 20128
rect 1336 20128 2536 20134
rect 1336 20125 1342 20128
rect 1422 20018 1428 20021
rect 228 20012 1428 20018
rect 2496 20018 2502 20021
rect 2496 20012 2536 20018
rect 228 19978 240 20012
rect 2524 19978 2536 20012
rect 228 19972 1428 19978
rect 1422 19969 1428 19972
rect 2496 19972 2536 19978
rect 2496 19969 2502 19972
rect 262 19862 268 19865
rect 228 19856 268 19862
rect 1336 19862 1342 19865
rect 1336 19856 2536 19862
rect 228 19822 240 19856
rect 2524 19822 2536 19856
rect 228 19816 268 19822
rect 262 19813 268 19816
rect 1336 19816 2536 19822
rect 1336 19813 1342 19816
rect 1422 19706 1428 19709
rect 228 19700 1428 19706
rect 2496 19706 2502 19709
rect 2496 19700 2536 19706
rect 228 19666 240 19700
rect 2524 19666 2536 19700
rect 228 19660 1428 19666
rect 1422 19657 1428 19660
rect 2496 19660 2536 19666
rect 2496 19657 2502 19660
rect 262 19550 268 19553
rect 228 19544 268 19550
rect 1336 19550 1342 19553
rect 1336 19544 2536 19550
rect 228 19510 240 19544
rect 2524 19510 2536 19544
rect 228 19504 268 19510
rect 262 19501 268 19504
rect 1336 19504 2536 19510
rect 1336 19501 1342 19504
rect 1422 19394 1428 19397
rect 228 19388 1428 19394
rect 2496 19394 2502 19397
rect 2496 19388 2536 19394
rect 228 19354 240 19388
rect 2524 19354 2536 19388
rect 228 19348 1428 19354
rect 1422 19345 1428 19348
rect 2496 19348 2536 19354
rect 2496 19345 2502 19348
rect 262 19238 268 19241
rect 228 19232 268 19238
rect 1336 19238 1342 19241
rect 1336 19232 2536 19238
rect 228 19198 240 19232
rect 2524 19198 2536 19232
rect 228 19192 268 19198
rect 262 19189 268 19192
rect 1336 19192 2536 19198
rect 1336 19189 1342 19192
rect 1422 19082 1428 19085
rect 228 19076 1428 19082
rect 2496 19082 2502 19085
rect 2496 19076 2536 19082
rect 228 19042 240 19076
rect 2524 19042 2536 19076
rect 228 19036 1428 19042
rect 1422 19033 1428 19036
rect 2496 19036 2536 19042
rect 2496 19033 2502 19036
rect 262 18926 268 18929
rect 228 18920 268 18926
rect 1336 18926 1342 18929
rect 1336 18920 2536 18926
rect 228 18886 240 18920
rect 2524 18886 2536 18920
rect 228 18880 268 18886
rect 262 18877 268 18880
rect 1336 18880 2536 18886
rect 1336 18877 1342 18880
rect 1422 18770 1428 18773
rect 228 18764 1428 18770
rect 2496 18770 2502 18773
rect 2496 18764 2536 18770
rect 228 18730 240 18764
rect 2524 18730 2536 18764
rect 228 18724 1428 18730
rect 1422 18721 1428 18724
rect 2496 18724 2536 18730
rect 2496 18721 2502 18724
rect 262 18614 268 18617
rect 228 18608 268 18614
rect 1336 18614 1342 18617
rect 1336 18608 2536 18614
rect 228 18574 240 18608
rect 2524 18574 2536 18608
rect 228 18568 268 18574
rect 262 18565 268 18568
rect 1336 18568 2536 18574
rect 1336 18565 1342 18568
rect 1422 18458 1428 18461
rect 228 18452 1428 18458
rect 2496 18458 2502 18461
rect 2496 18452 2536 18458
rect 228 18418 240 18452
rect 2524 18418 2536 18452
rect 228 18412 1428 18418
rect 1422 18409 1428 18412
rect 2496 18412 2536 18418
rect 2496 18409 2502 18412
rect 262 18302 268 18305
rect 228 18296 268 18302
rect 1336 18302 1342 18305
rect 1336 18296 2536 18302
rect 228 18262 240 18296
rect 2524 18262 2536 18296
rect 228 18256 268 18262
rect 262 18253 268 18256
rect 1336 18256 2536 18262
rect 1336 18253 1342 18256
rect 1422 18146 1428 18149
rect 228 18140 1428 18146
rect 2496 18146 2502 18149
rect 2496 18140 2536 18146
rect 228 18106 240 18140
rect 2524 18106 2536 18140
rect 228 18100 1428 18106
rect 1422 18097 1428 18100
rect 2496 18100 2536 18106
rect 2496 18097 2502 18100
rect 262 17990 268 17993
rect 228 17984 268 17990
rect 1336 17990 1342 17993
rect 1336 17984 2536 17990
rect 228 17950 240 17984
rect 2524 17950 2536 17984
rect 228 17944 268 17950
rect 262 17941 268 17944
rect 1336 17944 2536 17950
rect 1336 17941 1342 17944
rect 1422 17834 1428 17837
rect 228 17828 1428 17834
rect 2496 17834 2502 17837
rect 2496 17828 2536 17834
rect 228 17794 240 17828
rect 2524 17794 2536 17828
rect 228 17788 1428 17794
rect 1422 17785 1428 17788
rect 2496 17788 2536 17794
rect 2496 17785 2502 17788
rect 262 17678 268 17681
rect 228 17672 268 17678
rect 1336 17678 1342 17681
rect 1336 17672 2536 17678
rect 228 17638 240 17672
rect 2524 17638 2536 17672
rect 228 17632 268 17638
rect 262 17629 268 17632
rect 1336 17632 2536 17638
rect 1336 17629 1342 17632
rect 1422 17522 1428 17525
rect 228 17516 1428 17522
rect 2496 17522 2502 17525
rect 2496 17516 2536 17522
rect 228 17482 240 17516
rect 2524 17482 2536 17516
rect 228 17476 1428 17482
rect 1422 17473 1428 17476
rect 2496 17476 2536 17482
rect 2496 17473 2502 17476
rect 262 17366 268 17369
rect 228 17360 268 17366
rect 1336 17366 1342 17369
rect 1336 17360 2536 17366
rect 228 17326 240 17360
rect 2524 17326 2536 17360
rect 228 17320 268 17326
rect 262 17317 268 17320
rect 1336 17320 2536 17326
rect 1336 17317 1342 17320
rect 1422 17210 1428 17213
rect 228 17204 1428 17210
rect 2496 17210 2502 17213
rect 2496 17204 2536 17210
rect 228 17170 240 17204
rect 2524 17170 2536 17204
rect 228 17164 1428 17170
rect 1422 17161 1428 17164
rect 2496 17164 2536 17170
rect 2496 17161 2502 17164
rect 262 17054 268 17057
rect 228 17048 268 17054
rect 1336 17054 1342 17057
rect 1336 17048 2536 17054
rect 228 17014 240 17048
rect 2524 17014 2536 17048
rect 228 17008 268 17014
rect 262 17005 268 17008
rect 1336 17008 2536 17014
rect 1336 17005 1342 17008
rect 1422 16898 1428 16901
rect 228 16892 1428 16898
rect 2496 16898 2502 16901
rect 2496 16892 2536 16898
rect 228 16858 240 16892
rect 2524 16858 2536 16892
rect 228 16852 1428 16858
rect 1422 16849 1428 16852
rect 2496 16852 2536 16858
rect 2496 16849 2502 16852
rect 262 16742 268 16745
rect 228 16736 268 16742
rect 1336 16742 1342 16745
rect 1336 16736 2536 16742
rect 228 16702 240 16736
rect 2524 16702 2536 16736
rect 228 16696 268 16702
rect 262 16693 268 16696
rect 1336 16696 2536 16702
rect 1336 16693 1342 16696
rect 1422 16586 1428 16589
rect 228 16580 1428 16586
rect 2496 16586 2502 16589
rect 2496 16580 2536 16586
rect 228 16546 240 16580
rect 2524 16546 2536 16580
rect 228 16540 1428 16546
rect 1422 16537 1428 16540
rect 2496 16540 2536 16546
rect 2496 16537 2502 16540
rect 262 16430 268 16433
rect 228 16424 268 16430
rect 1336 16430 1342 16433
rect 1336 16424 2536 16430
rect 228 16390 240 16424
rect 2524 16390 2536 16424
rect 228 16384 268 16390
rect 262 16381 268 16384
rect 1336 16384 2536 16390
rect 1336 16381 1342 16384
rect 1422 16274 1428 16277
rect 228 16268 1428 16274
rect 2496 16274 2502 16277
rect 2496 16268 2536 16274
rect 228 16234 240 16268
rect 2524 16234 2536 16268
rect 228 16228 1428 16234
rect 1422 16225 1428 16228
rect 2496 16228 2536 16234
rect 2496 16225 2502 16228
rect 262 16118 268 16121
rect 228 16112 268 16118
rect 1336 16118 1342 16121
rect 1336 16112 2536 16118
rect 228 16078 240 16112
rect 2524 16078 2536 16112
rect 228 16072 268 16078
rect 262 16069 268 16072
rect 1336 16072 2536 16078
rect 1336 16069 1342 16072
rect 1422 15962 1428 15965
rect 228 15956 1428 15962
rect 2496 15962 2502 15965
rect 2496 15956 2536 15962
rect 228 15922 240 15956
rect 2524 15922 2536 15956
rect 228 15916 1428 15922
rect 1422 15913 1428 15916
rect 2496 15916 2536 15922
rect 2496 15913 2502 15916
rect 262 15806 268 15809
rect 228 15800 268 15806
rect 1336 15806 1342 15809
rect 1336 15800 2536 15806
rect 228 15766 240 15800
rect 2524 15766 2536 15800
rect 228 15760 268 15766
rect 262 15757 268 15760
rect 1336 15760 2536 15766
rect 1336 15757 1342 15760
rect 1422 15650 1428 15653
rect 228 15644 1428 15650
rect 2496 15650 2502 15653
rect 2496 15644 2536 15650
rect 228 15610 240 15644
rect 2524 15610 2536 15644
rect 228 15604 1428 15610
rect 1422 15601 1428 15604
rect 2496 15604 2536 15610
rect 2496 15601 2502 15604
rect 262 15494 268 15497
rect 228 15488 268 15494
rect 1336 15494 1342 15497
rect 1336 15488 2536 15494
rect 228 15454 240 15488
rect 2524 15454 2536 15488
rect 228 15448 268 15454
rect 262 15445 268 15448
rect 1336 15448 2536 15454
rect 1336 15445 1342 15448
rect 1422 15338 1428 15341
rect 228 15332 1428 15338
rect 2496 15338 2502 15341
rect 2496 15332 2536 15338
rect 228 15298 240 15332
rect 2524 15298 2536 15332
rect 228 15292 1428 15298
rect 1422 15289 1428 15292
rect 2496 15292 2536 15298
rect 2496 15289 2502 15292
rect 262 15182 268 15185
rect 228 15176 268 15182
rect 1336 15182 1342 15185
rect 1336 15176 2536 15182
rect 228 15142 240 15176
rect 2524 15142 2536 15176
rect 228 15136 268 15142
rect 262 15133 268 15136
rect 1336 15136 2536 15142
rect 1336 15133 1342 15136
rect 1422 15026 1428 15029
rect 228 15020 1428 15026
rect 2496 15026 2502 15029
rect 2496 15020 2536 15026
rect 228 14986 240 15020
rect 2524 14986 2536 15020
rect 228 14980 1428 14986
rect 1422 14977 1428 14980
rect 2496 14980 2536 14986
rect 2496 14977 2502 14980
rect 262 14870 268 14873
rect 228 14864 268 14870
rect 1336 14870 1342 14873
rect 1336 14864 2536 14870
rect 228 14830 240 14864
rect 2524 14830 2536 14864
rect 228 14824 268 14830
rect 262 14821 268 14824
rect 1336 14824 2536 14830
rect 1336 14821 1342 14824
rect 1422 14714 1428 14717
rect 228 14708 1428 14714
rect 2496 14714 2502 14717
rect 2496 14708 2536 14714
rect 228 14674 240 14708
rect 2524 14674 2536 14708
rect 228 14668 1428 14674
rect 1422 14665 1428 14668
rect 2496 14668 2536 14674
rect 2496 14665 2502 14668
rect 262 14558 268 14561
rect 228 14552 268 14558
rect 1336 14558 1342 14561
rect 1336 14552 2536 14558
rect 228 14518 240 14552
rect 2524 14518 2536 14552
rect 228 14512 268 14518
rect 262 14509 268 14512
rect 1336 14512 2536 14518
rect 1336 14509 1342 14512
rect 1422 14402 1428 14405
rect 228 14396 1428 14402
rect 2496 14402 2502 14405
rect 2496 14396 2536 14402
rect 228 14362 240 14396
rect 2524 14362 2536 14396
rect 228 14356 1428 14362
rect 1422 14353 1428 14356
rect 2496 14356 2536 14362
rect 2496 14353 2502 14356
rect 262 14246 268 14249
rect 228 14240 268 14246
rect 1336 14246 1342 14249
rect 1336 14240 2536 14246
rect 228 14206 240 14240
rect 2524 14206 2536 14240
rect 228 14200 268 14206
rect 262 14197 268 14200
rect 1336 14200 2536 14206
rect 1336 14197 1342 14200
rect 1422 14090 1428 14093
rect 228 14084 1428 14090
rect 2496 14090 2502 14093
rect 2496 14084 2536 14090
rect 228 14050 240 14084
rect 2524 14050 2536 14084
rect 228 14044 1428 14050
rect 1422 14041 1428 14044
rect 2496 14044 2536 14050
rect 2496 14041 2502 14044
rect 262 13934 268 13937
rect 228 13928 268 13934
rect 1336 13934 1342 13937
rect 1336 13928 2536 13934
rect 228 13894 240 13928
rect 2524 13894 2536 13928
rect 228 13888 268 13894
rect 262 13885 268 13888
rect 1336 13888 2536 13894
rect 1336 13885 1342 13888
rect 1422 13778 1428 13781
rect 228 13772 1428 13778
rect 2496 13778 2502 13781
rect 2496 13772 2536 13778
rect 228 13738 240 13772
rect 2524 13738 2536 13772
rect 228 13732 1428 13738
rect 1422 13729 1428 13732
rect 2496 13732 2536 13738
rect 2496 13729 2502 13732
rect 262 13622 268 13625
rect 228 13616 268 13622
rect 1336 13622 1342 13625
rect 1336 13616 2536 13622
rect 228 13582 240 13616
rect 2524 13582 2536 13616
rect 228 13576 268 13582
rect 262 13573 268 13576
rect 1336 13576 2536 13582
rect 1336 13573 1342 13576
rect 1422 13466 1428 13469
rect 228 13460 1428 13466
rect 2496 13466 2502 13469
rect 2496 13460 2536 13466
rect 228 13426 240 13460
rect 2524 13426 2536 13460
rect 228 13420 1428 13426
rect 1422 13417 1428 13420
rect 2496 13420 2536 13426
rect 2496 13417 2502 13420
rect 262 13310 268 13313
rect 228 13304 268 13310
rect 1336 13310 1342 13313
rect 1336 13304 2536 13310
rect 228 13270 240 13304
rect 2524 13270 2536 13304
rect 228 13264 268 13270
rect 262 13261 268 13264
rect 1336 13264 2536 13270
rect 1336 13261 1342 13264
rect 1422 13154 1428 13157
rect 228 13148 1428 13154
rect 2496 13154 2502 13157
rect 2496 13148 2536 13154
rect 228 13114 240 13148
rect 2524 13114 2536 13148
rect 228 13108 1428 13114
rect 1422 13105 1428 13108
rect 2496 13108 2536 13114
rect 2496 13105 2502 13108
rect 262 12998 268 13001
rect 228 12992 268 12998
rect 1336 12998 1342 13001
rect 1336 12992 2536 12998
rect 228 12958 240 12992
rect 2524 12958 2536 12992
rect 228 12952 268 12958
rect 262 12949 268 12952
rect 1336 12952 2536 12958
rect 1336 12949 1342 12952
rect 1422 12842 1428 12845
rect 228 12836 1428 12842
rect 2496 12842 2502 12845
rect 2496 12836 2536 12842
rect 228 12802 240 12836
rect 2524 12802 2536 12836
rect 228 12796 1428 12802
rect 1422 12793 1428 12796
rect 2496 12796 2536 12802
rect 2496 12793 2502 12796
rect 262 12686 268 12689
rect 228 12680 268 12686
rect 1336 12686 1342 12689
rect 1336 12680 2536 12686
rect 228 12646 240 12680
rect 2524 12646 2536 12680
rect 228 12640 268 12646
rect 262 12637 268 12640
rect 1336 12640 2536 12646
rect 1336 12637 1342 12640
rect 1422 12530 1428 12533
rect 228 12524 1428 12530
rect 2496 12530 2502 12533
rect 2496 12524 2536 12530
rect 228 12490 240 12524
rect 2524 12490 2536 12524
rect 228 12484 1428 12490
rect 1422 12481 1428 12484
rect 2496 12484 2536 12490
rect 2496 12481 2502 12484
rect 262 12374 268 12377
rect 228 12368 268 12374
rect 1336 12374 1342 12377
rect 1336 12368 2536 12374
rect 228 12334 240 12368
rect 2524 12334 2536 12368
rect 228 12328 268 12334
rect 262 12325 268 12328
rect 1336 12328 2536 12334
rect 1336 12325 1342 12328
rect 1422 12218 1428 12221
rect 228 12212 1428 12218
rect 2496 12218 2502 12221
rect 2496 12212 2536 12218
rect 228 12178 240 12212
rect 2524 12178 2536 12212
rect 228 12172 1428 12178
rect 1422 12169 1428 12172
rect 2496 12172 2536 12178
rect 2496 12169 2502 12172
rect 262 12062 268 12065
rect 228 12056 268 12062
rect 1336 12062 1342 12065
rect 1336 12056 2536 12062
rect 228 12022 240 12056
rect 2524 12022 2536 12056
rect 228 12016 268 12022
rect 262 12013 268 12016
rect 1336 12016 2536 12022
rect 1336 12013 1342 12016
rect 1422 11906 1428 11909
rect 228 11900 1428 11906
rect 2496 11906 2502 11909
rect 2496 11900 2536 11906
rect 228 11866 240 11900
rect 2524 11866 2536 11900
rect 228 11860 1428 11866
rect 1422 11857 1428 11860
rect 2496 11860 2536 11866
rect 2496 11857 2502 11860
rect 262 11750 268 11753
rect 228 11744 268 11750
rect 1336 11750 1342 11753
rect 1336 11744 2536 11750
rect 228 11710 240 11744
rect 2524 11710 2536 11744
rect 228 11704 268 11710
rect 262 11701 268 11704
rect 1336 11704 2536 11710
rect 1336 11701 1342 11704
rect 1422 11594 1428 11597
rect 228 11588 1428 11594
rect 2496 11594 2502 11597
rect 2496 11588 2536 11594
rect 228 11554 240 11588
rect 2524 11554 2536 11588
rect 228 11548 1428 11554
rect 1422 11545 1428 11548
rect 2496 11548 2536 11554
rect 2496 11545 2502 11548
rect 262 11438 268 11441
rect 228 11432 268 11438
rect 1336 11438 1342 11441
rect 1336 11432 2536 11438
rect 228 11398 240 11432
rect 2524 11398 2536 11432
rect 228 11392 268 11398
rect 262 11389 268 11392
rect 1336 11392 2536 11398
rect 1336 11389 1342 11392
rect 1422 11282 1428 11285
rect 228 11276 1428 11282
rect 2496 11282 2502 11285
rect 2496 11276 2536 11282
rect 228 11242 240 11276
rect 2524 11242 2536 11276
rect 228 11236 1428 11242
rect 1422 11233 1428 11236
rect 2496 11236 2536 11242
rect 2496 11233 2502 11236
rect 262 11126 268 11129
rect 228 11120 268 11126
rect 1336 11126 1342 11129
rect 1336 11120 2536 11126
rect 228 11086 240 11120
rect 2524 11086 2536 11120
rect 228 11080 268 11086
rect 262 11077 268 11080
rect 1336 11080 2536 11086
rect 1336 11077 1342 11080
rect 1422 10970 1428 10973
rect 228 10964 1428 10970
rect 2496 10970 2502 10973
rect 2496 10964 2536 10970
rect 228 10930 240 10964
rect 2524 10930 2536 10964
rect 228 10924 1428 10930
rect 1422 10921 1428 10924
rect 2496 10924 2536 10930
rect 2496 10921 2502 10924
rect 262 10814 268 10817
rect 228 10808 268 10814
rect 1336 10814 1342 10817
rect 1336 10808 2536 10814
rect 228 10774 240 10808
rect 2524 10774 2536 10808
rect 228 10768 268 10774
rect 262 10765 268 10768
rect 1336 10768 2536 10774
rect 1336 10765 1342 10768
rect 1422 10658 1428 10661
rect 228 10652 1428 10658
rect 2496 10658 2502 10661
rect 2496 10652 2536 10658
rect 228 10618 240 10652
rect 2524 10618 2536 10652
rect 228 10612 1428 10618
rect 1422 10609 1428 10612
rect 2496 10612 2536 10618
rect 2496 10609 2502 10612
rect 262 10502 268 10505
rect 228 10496 268 10502
rect 1336 10502 1342 10505
rect 1336 10496 2536 10502
rect 228 10462 240 10496
rect 2524 10462 2536 10496
rect 228 10456 268 10462
rect 262 10453 268 10456
rect 1336 10456 2536 10462
rect 1336 10453 1342 10456
rect 1422 10346 1428 10349
rect 228 10340 1428 10346
rect 2496 10346 2502 10349
rect 2496 10340 2536 10346
rect 228 10306 240 10340
rect 2524 10306 2536 10340
rect 228 10300 1428 10306
rect 1422 10297 1428 10300
rect 2496 10300 2536 10306
rect 2496 10297 2502 10300
rect 262 10190 268 10193
rect 228 10184 268 10190
rect 1336 10190 1342 10193
rect 1336 10184 2536 10190
rect 228 10150 240 10184
rect 2524 10150 2536 10184
rect 228 10144 268 10150
rect 262 10141 268 10144
rect 1336 10144 2536 10150
rect 1336 10141 1342 10144
rect 1422 10034 1428 10037
rect 228 10028 1428 10034
rect 2496 10034 2502 10037
rect 2496 10028 2536 10034
rect 228 9994 240 10028
rect 2524 9994 2536 10028
rect 228 9988 1428 9994
rect 1422 9985 1428 9988
rect 2496 9988 2536 9994
rect 2496 9985 2502 9988
rect 262 9878 268 9881
rect 228 9872 268 9878
rect 1336 9878 1342 9881
rect 1336 9872 2536 9878
rect 228 9838 240 9872
rect 2524 9838 2536 9872
rect 228 9832 268 9838
rect 262 9829 268 9832
rect 1336 9832 2536 9838
rect 1336 9829 1342 9832
rect 1422 9722 1428 9725
rect 228 9716 1428 9722
rect 2496 9722 2502 9725
rect 2496 9716 2536 9722
rect 228 9682 240 9716
rect 2524 9682 2536 9716
rect 228 9676 1428 9682
rect 1422 9673 1428 9676
rect 2496 9676 2536 9682
rect 2496 9673 2502 9676
rect 262 9566 268 9569
rect 228 9560 268 9566
rect 1336 9566 1342 9569
rect 1336 9560 2536 9566
rect 228 9526 240 9560
rect 2524 9526 2536 9560
rect 228 9520 268 9526
rect 262 9517 268 9520
rect 1336 9520 2536 9526
rect 1336 9517 1342 9520
rect 1422 9410 1428 9413
rect 228 9404 1428 9410
rect 2496 9410 2502 9413
rect 2496 9404 2536 9410
rect 228 9370 240 9404
rect 2524 9370 2536 9404
rect 228 9364 1428 9370
rect 1422 9361 1428 9364
rect 2496 9364 2536 9370
rect 2496 9361 2502 9364
rect 262 9254 268 9257
rect 228 9248 268 9254
rect 1336 9254 1342 9257
rect 1336 9248 2536 9254
rect 228 9214 240 9248
rect 2524 9214 2536 9248
rect 228 9208 268 9214
rect 262 9205 268 9208
rect 1336 9208 2536 9214
rect 1336 9205 1342 9208
rect 1422 9098 1428 9101
rect 228 9092 1428 9098
rect 2496 9098 2502 9101
rect 2496 9092 2536 9098
rect 228 9058 240 9092
rect 2524 9058 2536 9092
rect 228 9052 1428 9058
rect 1422 9049 1428 9052
rect 2496 9052 2536 9058
rect 2496 9049 2502 9052
rect 262 8942 268 8945
rect 228 8936 268 8942
rect 1336 8942 1342 8945
rect 1336 8936 2536 8942
rect 228 8902 240 8936
rect 2524 8902 2536 8936
rect 228 8896 268 8902
rect 262 8893 268 8896
rect 1336 8896 2536 8902
rect 1336 8893 1342 8896
rect 1422 8786 1428 8789
rect 228 8780 1428 8786
rect 2496 8786 2502 8789
rect 2496 8780 2536 8786
rect 228 8746 240 8780
rect 2524 8746 2536 8780
rect 228 8740 1428 8746
rect 1422 8737 1428 8740
rect 2496 8740 2536 8746
rect 2496 8737 2502 8740
rect 262 8630 268 8633
rect 228 8624 268 8630
rect 1336 8630 1342 8633
rect 1336 8624 2536 8630
rect 228 8590 240 8624
rect 2524 8590 2536 8624
rect 228 8584 268 8590
rect 262 8581 268 8584
rect 1336 8584 2536 8590
rect 1336 8581 1342 8584
rect 1422 8474 1428 8477
rect 228 8468 1428 8474
rect 2496 8474 2502 8477
rect 2496 8468 2536 8474
rect 228 8434 240 8468
rect 2524 8434 2536 8468
rect 228 8428 1428 8434
rect 1422 8425 1428 8428
rect 2496 8428 2536 8434
rect 2496 8425 2502 8428
rect 262 8318 268 8321
rect 228 8312 268 8318
rect 1336 8318 1342 8321
rect 1336 8312 2536 8318
rect 228 8278 240 8312
rect 2524 8278 2536 8312
rect 228 8272 268 8278
rect 262 8269 268 8272
rect 1336 8272 2536 8278
rect 1336 8269 1342 8272
rect 1422 8162 1428 8165
rect 228 8156 1428 8162
rect 2496 8162 2502 8165
rect 2496 8156 2536 8162
rect 228 8122 240 8156
rect 2524 8122 2536 8156
rect 228 8116 1428 8122
rect 1422 8113 1428 8116
rect 2496 8116 2536 8122
rect 2496 8113 2502 8116
rect 262 8006 268 8009
rect 228 8000 268 8006
rect 1336 8006 1342 8009
rect 1336 8000 2536 8006
rect 228 7966 240 8000
rect 2524 7966 2536 8000
rect 228 7960 268 7966
rect 262 7957 268 7960
rect 1336 7960 2536 7966
rect 1336 7957 1342 7960
rect 1422 7850 1428 7853
rect 228 7844 1428 7850
rect 2496 7850 2502 7853
rect 2496 7844 2536 7850
rect 228 7810 240 7844
rect 2524 7810 2536 7844
rect 228 7804 1428 7810
rect 1422 7801 1428 7804
rect 2496 7804 2536 7810
rect 2496 7801 2502 7804
rect 262 7694 268 7697
rect 228 7688 268 7694
rect 1336 7694 1342 7697
rect 1336 7688 2536 7694
rect 228 7654 240 7688
rect 2524 7654 2536 7688
rect 228 7648 268 7654
rect 262 7645 268 7648
rect 1336 7648 2536 7654
rect 1336 7645 1342 7648
rect 1422 7538 1428 7541
rect 228 7532 1428 7538
rect 2496 7538 2502 7541
rect 2496 7532 2536 7538
rect 228 7498 240 7532
rect 2524 7498 2536 7532
rect 228 7492 1428 7498
rect 1422 7489 1428 7492
rect 2496 7492 2536 7498
rect 2496 7489 2502 7492
rect 262 7382 268 7385
rect 228 7376 268 7382
rect 1336 7382 1342 7385
rect 1336 7376 2536 7382
rect 228 7342 240 7376
rect 2524 7342 2536 7376
rect 228 7336 268 7342
rect 262 7333 268 7336
rect 1336 7336 2536 7342
rect 1336 7333 1342 7336
rect 1422 7226 1428 7229
rect 228 7220 1428 7226
rect 2496 7226 2502 7229
rect 2496 7220 2536 7226
rect 228 7186 240 7220
rect 2524 7186 2536 7220
rect 228 7180 1428 7186
rect 1422 7177 1428 7180
rect 2496 7180 2536 7186
rect 2496 7177 2502 7180
rect 262 7070 268 7073
rect 228 7064 268 7070
rect 1336 7070 1342 7073
rect 1336 7064 2536 7070
rect 228 7030 240 7064
rect 2524 7030 2536 7064
rect 228 7024 268 7030
rect 262 7021 268 7024
rect 1336 7024 2536 7030
rect 1336 7021 1342 7024
rect 1422 6914 1428 6917
rect 228 6908 1428 6914
rect 2496 6914 2502 6917
rect 2496 6908 2536 6914
rect 228 6874 240 6908
rect 2524 6874 2536 6908
rect 228 6868 1428 6874
rect 1422 6865 1428 6868
rect 2496 6868 2536 6874
rect 2496 6865 2502 6868
rect 262 6758 268 6761
rect 228 6752 268 6758
rect 1336 6758 1342 6761
rect 1336 6752 2536 6758
rect 228 6718 240 6752
rect 2524 6718 2536 6752
rect 228 6712 268 6718
rect 262 6709 268 6712
rect 1336 6712 2536 6718
rect 1336 6709 1342 6712
rect 1422 6602 1428 6605
rect 228 6596 1428 6602
rect 2496 6602 2502 6605
rect 2496 6596 2536 6602
rect 228 6562 240 6596
rect 2524 6562 2536 6596
rect 228 6556 1428 6562
rect 1422 6553 1428 6556
rect 2496 6556 2536 6562
rect 2496 6553 2502 6556
rect 262 6446 268 6449
rect 228 6440 268 6446
rect 1336 6446 1342 6449
rect 1336 6440 2536 6446
rect 228 6406 240 6440
rect 2524 6406 2536 6440
rect 228 6400 268 6406
rect 262 6397 268 6400
rect 1336 6400 2536 6406
rect 1336 6397 1342 6400
rect 1422 6290 1428 6293
rect 228 6284 1428 6290
rect 2496 6290 2502 6293
rect 2496 6284 2536 6290
rect 228 6250 240 6284
rect 2524 6250 2536 6284
rect 228 6244 1428 6250
rect 1422 6241 1428 6244
rect 2496 6244 2536 6250
rect 2496 6241 2502 6244
rect 262 6134 268 6137
rect 228 6128 268 6134
rect 1336 6134 1342 6137
rect 1336 6128 2536 6134
rect 228 6094 240 6128
rect 2524 6094 2536 6128
rect 228 6088 268 6094
rect 262 6085 268 6088
rect 1336 6088 2536 6094
rect 1336 6085 1342 6088
rect 1422 5978 1428 5981
rect 228 5972 1428 5978
rect 2496 5978 2502 5981
rect 2496 5972 2536 5978
rect 228 5938 240 5972
rect 2524 5938 2536 5972
rect 228 5932 1428 5938
rect 1422 5929 1428 5932
rect 2496 5932 2536 5938
rect 2496 5929 2502 5932
rect 262 5822 268 5825
rect 228 5816 268 5822
rect 1336 5822 1342 5825
rect 1336 5816 2536 5822
rect 228 5782 240 5816
rect 2524 5782 2536 5816
rect 228 5776 268 5782
rect 262 5773 268 5776
rect 1336 5776 2536 5782
rect 1336 5773 1342 5776
rect 1422 5666 1428 5669
rect 228 5660 1428 5666
rect 2496 5666 2502 5669
rect 2496 5660 2536 5666
rect 228 5626 240 5660
rect 2524 5626 2536 5660
rect 228 5620 1428 5626
rect 1422 5617 1428 5620
rect 2496 5620 2536 5626
rect 2496 5617 2502 5620
rect 262 5510 268 5513
rect 228 5504 268 5510
rect 1336 5510 1342 5513
rect 1336 5504 2536 5510
rect 228 5470 240 5504
rect 2524 5470 2536 5504
rect 228 5464 268 5470
rect 262 5461 268 5464
rect 1336 5464 2536 5470
rect 1336 5461 1342 5464
rect 1422 5354 1428 5357
rect 228 5348 1428 5354
rect 2496 5354 2502 5357
rect 2496 5348 2536 5354
rect 228 5314 240 5348
rect 2524 5314 2536 5348
rect 228 5308 1428 5314
rect 1422 5305 1428 5308
rect 2496 5308 2536 5314
rect 2496 5305 2502 5308
rect 262 5198 268 5201
rect 228 5192 268 5198
rect 1336 5198 1342 5201
rect 1336 5192 2536 5198
rect 228 5158 240 5192
rect 2524 5158 2536 5192
rect 228 5152 268 5158
rect 262 5149 268 5152
rect 1336 5152 2536 5158
rect 1336 5149 1342 5152
rect 1422 5042 1428 5045
rect 228 5036 1428 5042
rect 2496 5042 2502 5045
rect 2496 5036 2536 5042
rect 228 5002 240 5036
rect 2524 5002 2536 5036
rect 228 4996 1428 5002
rect 1422 4993 1428 4996
rect 2496 4996 2536 5002
rect 2496 4993 2502 4996
rect 262 4886 268 4889
rect 228 4880 268 4886
rect 1336 4886 1342 4889
rect 1336 4880 2536 4886
rect 228 4846 240 4880
rect 2524 4846 2536 4880
rect 228 4840 268 4846
rect 262 4837 268 4840
rect 1336 4840 2536 4846
rect 1336 4837 1342 4840
rect 1422 4730 1428 4733
rect 228 4724 1428 4730
rect 2496 4730 2502 4733
rect 2496 4724 2536 4730
rect 228 4690 240 4724
rect 2524 4690 2536 4724
rect 228 4684 1428 4690
rect 1422 4681 1428 4684
rect 2496 4684 2536 4690
rect 2496 4681 2502 4684
rect 262 4574 268 4577
rect 228 4568 268 4574
rect 1336 4574 1342 4577
rect 1336 4568 2536 4574
rect 228 4534 240 4568
rect 2524 4534 2536 4568
rect 228 4528 268 4534
rect 262 4525 268 4528
rect 1336 4528 2536 4534
rect 1336 4525 1342 4528
rect 1422 4418 1428 4421
rect 228 4412 1428 4418
rect 2496 4418 2502 4421
rect 2496 4412 2536 4418
rect 228 4378 240 4412
rect 2524 4378 2536 4412
rect 228 4372 1428 4378
rect 1422 4369 1428 4372
rect 2496 4372 2536 4378
rect 2496 4369 2502 4372
rect 262 4262 268 4265
rect 228 4256 268 4262
rect 1336 4262 1342 4265
rect 1336 4256 2536 4262
rect 228 4222 240 4256
rect 2524 4222 2536 4256
rect 228 4216 268 4222
rect 262 4213 268 4216
rect 1336 4216 2536 4222
rect 1336 4213 1342 4216
rect 1422 4106 1428 4109
rect 228 4100 1428 4106
rect 2496 4106 2502 4109
rect 2496 4100 2536 4106
rect 228 4066 240 4100
rect 2524 4066 2536 4100
rect 228 4060 1428 4066
rect 1422 4057 1428 4060
rect 2496 4060 2536 4066
rect 2496 4057 2502 4060
rect 262 3950 268 3953
rect 228 3944 268 3950
rect 1336 3950 1342 3953
rect 1336 3944 2536 3950
rect 228 3910 240 3944
rect 2524 3910 2536 3944
rect 228 3904 268 3910
rect 262 3901 268 3904
rect 1336 3904 2536 3910
rect 1336 3901 1342 3904
rect 1422 3794 1428 3797
rect 228 3788 1428 3794
rect 2496 3794 2502 3797
rect 2496 3788 2536 3794
rect 228 3754 240 3788
rect 2524 3754 2536 3788
rect 228 3748 1428 3754
rect 1422 3745 1428 3748
rect 2496 3748 2536 3754
rect 2496 3745 2502 3748
rect 262 3638 268 3641
rect 228 3632 268 3638
rect 1336 3638 1342 3641
rect 1336 3632 2536 3638
rect 228 3598 240 3632
rect 2524 3598 2536 3632
rect 228 3592 268 3598
rect 262 3589 268 3592
rect 1336 3592 2536 3598
rect 1336 3589 1342 3592
rect 1422 3482 1428 3485
rect 228 3476 1428 3482
rect 2496 3482 2502 3485
rect 2496 3476 2536 3482
rect 228 3442 240 3476
rect 2524 3442 2536 3476
rect 228 3436 1428 3442
rect 1422 3433 1428 3436
rect 2496 3436 2536 3442
rect 2496 3433 2502 3436
rect 262 3326 268 3329
rect 228 3320 268 3326
rect 1336 3326 1342 3329
rect 1336 3320 2536 3326
rect 228 3286 240 3320
rect 2524 3286 2536 3320
rect 228 3280 268 3286
rect 262 3277 268 3280
rect 1336 3280 2536 3286
rect 1336 3277 1342 3280
rect 1422 3170 1428 3173
rect 228 3164 1428 3170
rect 2496 3170 2502 3173
rect 2496 3164 2536 3170
rect 228 3130 240 3164
rect 2524 3130 2536 3164
rect 228 3124 1428 3130
rect 1422 3121 1428 3124
rect 2496 3124 2536 3130
rect 2496 3121 2502 3124
rect 262 3014 268 3017
rect 228 3008 268 3014
rect 1336 3014 1342 3017
rect 1336 3008 2536 3014
rect 228 2974 240 3008
rect 2524 2974 2536 3008
rect 228 2968 268 2974
rect 262 2965 268 2968
rect 1336 2968 2536 2974
rect 1336 2965 1342 2968
rect 1422 2858 1428 2861
rect 228 2852 1428 2858
rect 2496 2858 2502 2861
rect 2496 2852 2536 2858
rect 228 2818 240 2852
rect 2524 2818 2536 2852
rect 228 2812 1428 2818
rect 1422 2809 1428 2812
rect 2496 2812 2536 2818
rect 2496 2809 2502 2812
rect 262 2702 268 2705
rect 228 2696 268 2702
rect 1336 2702 1342 2705
rect 1336 2696 2536 2702
rect 228 2662 240 2696
rect 2524 2662 2536 2696
rect 228 2656 268 2662
rect 262 2653 268 2656
rect 1336 2656 2536 2662
rect 1336 2653 1342 2656
rect 1422 2546 1428 2549
rect 228 2540 1428 2546
rect 2496 2546 2502 2549
rect 2496 2540 2536 2546
rect 228 2506 240 2540
rect 2524 2506 2536 2540
rect 228 2500 1428 2506
rect 1422 2497 1428 2500
rect 2496 2500 2536 2506
rect 2496 2497 2502 2500
rect 262 2390 268 2393
rect 228 2384 268 2390
rect 1336 2390 1342 2393
rect 1336 2384 2536 2390
rect 228 2350 240 2384
rect 2524 2350 2536 2384
rect 228 2344 268 2350
rect 262 2341 268 2344
rect 1336 2344 2536 2350
rect 1336 2341 1342 2344
rect 1422 2234 1428 2237
rect 228 2228 1428 2234
rect 2496 2234 2502 2237
rect 2496 2228 2536 2234
rect 228 2194 240 2228
rect 2524 2194 2536 2228
rect 228 2188 1428 2194
rect 1422 2185 1428 2188
rect 2496 2188 2536 2194
rect 2496 2185 2502 2188
rect 262 2078 268 2081
rect 228 2072 268 2078
rect 1336 2078 1342 2081
rect 1336 2072 2536 2078
rect 228 2038 240 2072
rect 2524 2038 2536 2072
rect 228 2032 268 2038
rect 262 2029 268 2032
rect 1336 2032 2536 2038
rect 1336 2029 1342 2032
rect 1422 1922 1428 1925
rect 228 1916 1428 1922
rect 2496 1922 2502 1925
rect 2496 1916 2536 1922
rect 228 1882 240 1916
rect 2524 1882 2536 1916
rect 228 1876 1428 1882
rect 1422 1873 1428 1876
rect 2496 1876 2536 1882
rect 2496 1873 2502 1876
rect 262 1766 268 1769
rect 228 1760 268 1766
rect 1336 1766 1342 1769
rect 1336 1760 2536 1766
rect 228 1726 240 1760
rect 2524 1726 2536 1760
rect 228 1720 268 1726
rect 262 1717 268 1720
rect 1336 1720 2536 1726
rect 1336 1717 1342 1720
rect 1422 1610 1428 1613
rect 228 1604 1428 1610
rect 2496 1610 2502 1613
rect 2496 1604 2536 1610
rect 228 1570 240 1604
rect 2524 1570 2536 1604
rect 228 1564 1428 1570
rect 1422 1561 1428 1564
rect 2496 1564 2536 1570
rect 2496 1561 2502 1564
rect 262 1454 268 1457
rect 228 1448 268 1454
rect 1336 1454 1342 1457
rect 1336 1448 2536 1454
rect 228 1414 240 1448
rect 2524 1414 2536 1448
rect 228 1408 268 1414
rect 262 1405 268 1408
rect 1336 1408 2536 1414
rect 1336 1405 1342 1408
rect 1422 1298 1428 1301
rect 228 1292 1428 1298
rect 2496 1298 2502 1301
rect 2496 1292 2536 1298
rect 228 1258 240 1292
rect 2524 1258 2536 1292
rect 228 1252 1428 1258
rect 1422 1249 1428 1252
rect 2496 1252 2536 1258
rect 2496 1249 2502 1252
rect 262 1142 268 1145
rect 228 1136 268 1142
rect 1336 1142 1342 1145
rect 1336 1136 2536 1142
rect 228 1102 240 1136
rect 2524 1102 2536 1136
rect 228 1096 268 1102
rect 262 1093 268 1096
rect 1336 1096 2536 1102
rect 1336 1093 1342 1096
rect 1422 986 1428 989
rect 228 980 1428 986
rect 2496 986 2502 989
rect 2496 980 2536 986
rect 228 946 240 980
rect 2524 946 2536 980
rect 228 940 1428 946
rect 1422 937 1428 940
rect 2496 940 2536 946
rect 2496 937 2502 940
rect 262 830 268 833
rect 228 824 268 830
rect 1336 830 1342 833
rect 1336 824 2536 830
rect 228 790 240 824
rect 2524 790 2536 824
rect 228 784 268 790
rect 262 781 268 784
rect 1336 784 2536 790
rect 1336 781 1342 784
rect 1422 674 1428 677
rect 228 668 1428 674
rect 2496 674 2502 677
rect 2496 668 2536 674
rect 228 634 240 668
rect 2524 634 2536 668
rect 228 628 1428 634
rect 1422 625 1428 628
rect 2496 628 2536 634
rect 2496 625 2502 628
rect 262 518 268 521
rect 228 512 268 518
rect 1336 518 1342 521
rect 1336 512 2536 518
rect 228 478 240 512
rect 2524 478 2536 512
rect 228 472 268 478
rect 262 469 268 472
rect 1336 472 2536 478
rect 1336 469 1342 472
rect 1422 362 1428 365
rect 228 356 1428 362
rect 2496 362 2502 365
rect 2496 356 2536 362
rect 228 322 240 356
rect 2524 322 2536 356
rect 228 316 1428 322
rect 1422 313 1428 316
rect 2496 316 2536 322
rect 2496 313 2502 316
rect 140 227 194 233
rect 262 206 268 209
rect 228 200 268 206
rect 1336 206 1342 209
rect 1336 200 2536 206
rect 228 166 240 200
rect 2524 166 2536 200
rect 228 160 268 166
rect 262 157 268 160
rect 1336 160 2536 166
rect 1336 157 1342 160
rect 60 106 106 130
rect 2580 130 2586 42980
rect 2620 130 2626 42980
rect 2580 106 2626 130
rect 60 100 2626 106
rect 60 66 130 100
rect 2556 66 2626 100
rect 60 60 2626 66
<< via1 >>
rect 268 42944 1336 42953
rect 268 42910 1336 42944
rect 268 42901 1336 42910
rect 140 42871 194 42877
rect 140 239 150 42871
rect 150 239 184 42871
rect 184 239 194 42871
rect 1428 42788 2496 42797
rect 1428 42754 2496 42788
rect 1428 42745 2496 42754
rect 268 42632 1336 42641
rect 268 42598 1336 42632
rect 268 42589 1336 42598
rect 1428 42476 2496 42485
rect 1428 42442 2496 42476
rect 1428 42433 2496 42442
rect 268 42320 1336 42329
rect 268 42286 1336 42320
rect 268 42277 1336 42286
rect 1428 42164 2496 42173
rect 1428 42130 2496 42164
rect 1428 42121 2496 42130
rect 268 42008 1336 42017
rect 268 41974 1336 42008
rect 268 41965 1336 41974
rect 1428 41852 2496 41861
rect 1428 41818 2496 41852
rect 1428 41809 2496 41818
rect 268 41696 1336 41705
rect 268 41662 1336 41696
rect 268 41653 1336 41662
rect 1428 41540 2496 41549
rect 1428 41506 2496 41540
rect 1428 41497 2496 41506
rect 268 41384 1336 41393
rect 268 41350 1336 41384
rect 268 41341 1336 41350
rect 1428 41228 2496 41237
rect 1428 41194 2496 41228
rect 1428 41185 2496 41194
rect 268 41072 1336 41081
rect 268 41038 1336 41072
rect 268 41029 1336 41038
rect 1428 40916 2496 40925
rect 1428 40882 2496 40916
rect 1428 40873 2496 40882
rect 268 40760 1336 40769
rect 268 40726 1336 40760
rect 268 40717 1336 40726
rect 1428 40604 2496 40613
rect 1428 40570 2496 40604
rect 1428 40561 2496 40570
rect 268 40448 1336 40457
rect 268 40414 1336 40448
rect 268 40405 1336 40414
rect 1428 40292 2496 40301
rect 1428 40258 2496 40292
rect 1428 40249 2496 40258
rect 268 40136 1336 40145
rect 268 40102 1336 40136
rect 268 40093 1336 40102
rect 1428 39980 2496 39989
rect 1428 39946 2496 39980
rect 1428 39937 2496 39946
rect 268 39824 1336 39833
rect 268 39790 1336 39824
rect 268 39781 1336 39790
rect 1428 39668 2496 39677
rect 1428 39634 2496 39668
rect 1428 39625 2496 39634
rect 268 39512 1336 39521
rect 268 39478 1336 39512
rect 268 39469 1336 39478
rect 1428 39356 2496 39365
rect 1428 39322 2496 39356
rect 1428 39313 2496 39322
rect 268 39200 1336 39209
rect 268 39166 1336 39200
rect 268 39157 1336 39166
rect 1428 39044 2496 39053
rect 1428 39010 2496 39044
rect 1428 39001 2496 39010
rect 268 38888 1336 38897
rect 268 38854 1336 38888
rect 268 38845 1336 38854
rect 1428 38732 2496 38741
rect 1428 38698 2496 38732
rect 1428 38689 2496 38698
rect 268 38576 1336 38585
rect 268 38542 1336 38576
rect 268 38533 1336 38542
rect 1428 38420 2496 38429
rect 1428 38386 2496 38420
rect 1428 38377 2496 38386
rect 268 38264 1336 38273
rect 268 38230 1336 38264
rect 268 38221 1336 38230
rect 1428 38108 2496 38117
rect 1428 38074 2496 38108
rect 1428 38065 2496 38074
rect 268 37952 1336 37961
rect 268 37918 1336 37952
rect 268 37909 1336 37918
rect 1428 37796 2496 37805
rect 1428 37762 2496 37796
rect 1428 37753 2496 37762
rect 268 37640 1336 37649
rect 268 37606 1336 37640
rect 268 37597 1336 37606
rect 1428 37484 2496 37493
rect 1428 37450 2496 37484
rect 1428 37441 2496 37450
rect 268 37328 1336 37337
rect 268 37294 1336 37328
rect 268 37285 1336 37294
rect 1428 37172 2496 37181
rect 1428 37138 2496 37172
rect 1428 37129 2496 37138
rect 268 37016 1336 37025
rect 268 36982 1336 37016
rect 268 36973 1336 36982
rect 1428 36860 2496 36869
rect 1428 36826 2496 36860
rect 1428 36817 2496 36826
rect 268 36704 1336 36713
rect 268 36670 1336 36704
rect 268 36661 1336 36670
rect 1428 36548 2496 36557
rect 1428 36514 2496 36548
rect 1428 36505 2496 36514
rect 268 36392 1336 36401
rect 268 36358 1336 36392
rect 268 36349 1336 36358
rect 1428 36236 2496 36245
rect 1428 36202 2496 36236
rect 1428 36193 2496 36202
rect 268 36080 1336 36089
rect 268 36046 1336 36080
rect 268 36037 1336 36046
rect 1428 35924 2496 35933
rect 1428 35890 2496 35924
rect 1428 35881 2496 35890
rect 268 35768 1336 35777
rect 268 35734 1336 35768
rect 268 35725 1336 35734
rect 1428 35612 2496 35621
rect 1428 35578 2496 35612
rect 1428 35569 2496 35578
rect 268 35456 1336 35465
rect 268 35422 1336 35456
rect 268 35413 1336 35422
rect 1428 35300 2496 35309
rect 1428 35266 2496 35300
rect 1428 35257 2496 35266
rect 268 35144 1336 35153
rect 268 35110 1336 35144
rect 268 35101 1336 35110
rect 1428 34988 2496 34997
rect 1428 34954 2496 34988
rect 1428 34945 2496 34954
rect 268 34832 1336 34841
rect 268 34798 1336 34832
rect 268 34789 1336 34798
rect 1428 34676 2496 34685
rect 1428 34642 2496 34676
rect 1428 34633 2496 34642
rect 268 34520 1336 34529
rect 268 34486 1336 34520
rect 268 34477 1336 34486
rect 1428 34364 2496 34373
rect 1428 34330 2496 34364
rect 1428 34321 2496 34330
rect 268 34208 1336 34217
rect 268 34174 1336 34208
rect 268 34165 1336 34174
rect 1428 34052 2496 34061
rect 1428 34018 2496 34052
rect 1428 34009 2496 34018
rect 268 33896 1336 33905
rect 268 33862 1336 33896
rect 268 33853 1336 33862
rect 1428 33740 2496 33749
rect 1428 33706 2496 33740
rect 1428 33697 2496 33706
rect 268 33584 1336 33593
rect 268 33550 1336 33584
rect 268 33541 1336 33550
rect 1428 33428 2496 33437
rect 1428 33394 2496 33428
rect 1428 33385 2496 33394
rect 268 33272 1336 33281
rect 268 33238 1336 33272
rect 268 33229 1336 33238
rect 1428 33116 2496 33125
rect 1428 33082 2496 33116
rect 1428 33073 2496 33082
rect 268 32960 1336 32969
rect 268 32926 1336 32960
rect 268 32917 1336 32926
rect 1428 32804 2496 32813
rect 1428 32770 2496 32804
rect 1428 32761 2496 32770
rect 268 32648 1336 32657
rect 268 32614 1336 32648
rect 268 32605 1336 32614
rect 1428 32492 2496 32501
rect 1428 32458 2496 32492
rect 1428 32449 2496 32458
rect 268 32336 1336 32345
rect 268 32302 1336 32336
rect 268 32293 1336 32302
rect 1428 32180 2496 32189
rect 1428 32146 2496 32180
rect 1428 32137 2496 32146
rect 268 32024 1336 32033
rect 268 31990 1336 32024
rect 268 31981 1336 31990
rect 1428 31868 2496 31877
rect 1428 31834 2496 31868
rect 1428 31825 2496 31834
rect 268 31712 1336 31721
rect 268 31678 1336 31712
rect 268 31669 1336 31678
rect 1428 31556 2496 31565
rect 1428 31522 2496 31556
rect 1428 31513 2496 31522
rect 268 31400 1336 31409
rect 268 31366 1336 31400
rect 268 31357 1336 31366
rect 1428 31244 2496 31253
rect 1428 31210 2496 31244
rect 1428 31201 2496 31210
rect 268 31088 1336 31097
rect 268 31054 1336 31088
rect 268 31045 1336 31054
rect 1428 30932 2496 30941
rect 1428 30898 2496 30932
rect 1428 30889 2496 30898
rect 268 30776 1336 30785
rect 268 30742 1336 30776
rect 268 30733 1336 30742
rect 1428 30620 2496 30629
rect 1428 30586 2496 30620
rect 1428 30577 2496 30586
rect 268 30464 1336 30473
rect 268 30430 1336 30464
rect 268 30421 1336 30430
rect 1428 30308 2496 30317
rect 1428 30274 2496 30308
rect 1428 30265 2496 30274
rect 268 30152 1336 30161
rect 268 30118 1336 30152
rect 268 30109 1336 30118
rect 1428 29996 2496 30005
rect 1428 29962 2496 29996
rect 1428 29953 2496 29962
rect 268 29840 1336 29849
rect 268 29806 1336 29840
rect 268 29797 1336 29806
rect 1428 29684 2496 29693
rect 1428 29650 2496 29684
rect 1428 29641 2496 29650
rect 268 29528 1336 29537
rect 268 29494 1336 29528
rect 268 29485 1336 29494
rect 1428 29372 2496 29381
rect 1428 29338 2496 29372
rect 1428 29329 2496 29338
rect 268 29216 1336 29225
rect 268 29182 1336 29216
rect 268 29173 1336 29182
rect 1428 29060 2496 29069
rect 1428 29026 2496 29060
rect 1428 29017 2496 29026
rect 268 28904 1336 28913
rect 268 28870 1336 28904
rect 268 28861 1336 28870
rect 1428 28748 2496 28757
rect 1428 28714 2496 28748
rect 1428 28705 2496 28714
rect 268 28592 1336 28601
rect 268 28558 1336 28592
rect 268 28549 1336 28558
rect 1428 28436 2496 28445
rect 1428 28402 2496 28436
rect 1428 28393 2496 28402
rect 268 28280 1336 28289
rect 268 28246 1336 28280
rect 268 28237 1336 28246
rect 1428 28124 2496 28133
rect 1428 28090 2496 28124
rect 1428 28081 2496 28090
rect 268 27968 1336 27977
rect 268 27934 1336 27968
rect 268 27925 1336 27934
rect 1428 27812 2496 27821
rect 1428 27778 2496 27812
rect 1428 27769 2496 27778
rect 268 27656 1336 27665
rect 268 27622 1336 27656
rect 268 27613 1336 27622
rect 1428 27500 2496 27509
rect 1428 27466 2496 27500
rect 1428 27457 2496 27466
rect 268 27344 1336 27353
rect 268 27310 1336 27344
rect 268 27301 1336 27310
rect 1428 27188 2496 27197
rect 1428 27154 2496 27188
rect 1428 27145 2496 27154
rect 268 27032 1336 27041
rect 268 26998 1336 27032
rect 268 26989 1336 26998
rect 1428 26876 2496 26885
rect 1428 26842 2496 26876
rect 1428 26833 2496 26842
rect 268 26720 1336 26729
rect 268 26686 1336 26720
rect 268 26677 1336 26686
rect 1428 26564 2496 26573
rect 1428 26530 2496 26564
rect 1428 26521 2496 26530
rect 268 26408 1336 26417
rect 268 26374 1336 26408
rect 268 26365 1336 26374
rect 1428 26252 2496 26261
rect 1428 26218 2496 26252
rect 1428 26209 2496 26218
rect 268 26096 1336 26105
rect 268 26062 1336 26096
rect 268 26053 1336 26062
rect 1428 25940 2496 25949
rect 1428 25906 2496 25940
rect 1428 25897 2496 25906
rect 268 25784 1336 25793
rect 268 25750 1336 25784
rect 268 25741 1336 25750
rect 1428 25628 2496 25637
rect 1428 25594 2496 25628
rect 1428 25585 2496 25594
rect 268 25472 1336 25481
rect 268 25438 1336 25472
rect 268 25429 1336 25438
rect 1428 25316 2496 25325
rect 1428 25282 2496 25316
rect 1428 25273 2496 25282
rect 268 25160 1336 25169
rect 268 25126 1336 25160
rect 268 25117 1336 25126
rect 1428 25004 2496 25013
rect 1428 24970 2496 25004
rect 1428 24961 2496 24970
rect 268 24848 1336 24857
rect 268 24814 1336 24848
rect 268 24805 1336 24814
rect 1428 24692 2496 24701
rect 1428 24658 2496 24692
rect 1428 24649 2496 24658
rect 268 24536 1336 24545
rect 268 24502 1336 24536
rect 268 24493 1336 24502
rect 1428 24380 2496 24389
rect 1428 24346 2496 24380
rect 1428 24337 2496 24346
rect 268 24224 1336 24233
rect 268 24190 1336 24224
rect 268 24181 1336 24190
rect 1428 24068 2496 24077
rect 1428 24034 2496 24068
rect 1428 24025 2496 24034
rect 268 23912 1336 23921
rect 268 23878 1336 23912
rect 268 23869 1336 23878
rect 1428 23756 2496 23765
rect 1428 23722 2496 23756
rect 1428 23713 2496 23722
rect 268 23600 1336 23609
rect 268 23566 1336 23600
rect 268 23557 1336 23566
rect 1428 23444 2496 23453
rect 1428 23410 2496 23444
rect 1428 23401 2496 23410
rect 268 23288 1336 23297
rect 268 23254 1336 23288
rect 268 23245 1336 23254
rect 1428 23132 2496 23141
rect 1428 23098 2496 23132
rect 1428 23089 2496 23098
rect 268 22976 1336 22985
rect 268 22942 1336 22976
rect 268 22933 1336 22942
rect 1428 22820 2496 22829
rect 1428 22786 2496 22820
rect 1428 22777 2496 22786
rect 268 22664 1336 22673
rect 268 22630 1336 22664
rect 268 22621 1336 22630
rect 1428 22508 2496 22517
rect 1428 22474 2496 22508
rect 1428 22465 2496 22474
rect 268 22352 1336 22361
rect 268 22318 1336 22352
rect 268 22309 1336 22318
rect 1428 22196 2496 22205
rect 1428 22162 2496 22196
rect 1428 22153 2496 22162
rect 268 22040 1336 22049
rect 268 22006 1336 22040
rect 268 21997 1336 22006
rect 1428 21884 2496 21893
rect 1428 21850 2496 21884
rect 1428 21841 2496 21850
rect 268 21728 1336 21737
rect 268 21694 1336 21728
rect 268 21685 1336 21694
rect 1428 21572 2496 21581
rect 1428 21538 2496 21572
rect 1428 21529 2496 21538
rect 268 21416 1336 21425
rect 268 21382 1336 21416
rect 268 21373 1336 21382
rect 1428 21260 2496 21269
rect 1428 21226 2496 21260
rect 1428 21217 2496 21226
rect 268 21104 1336 21113
rect 268 21070 1336 21104
rect 268 21061 1336 21070
rect 1428 20948 2496 20957
rect 1428 20914 2496 20948
rect 1428 20905 2496 20914
rect 268 20792 1336 20801
rect 268 20758 1336 20792
rect 268 20749 1336 20758
rect 1428 20636 2496 20645
rect 1428 20602 2496 20636
rect 1428 20593 2496 20602
rect 268 20480 1336 20489
rect 268 20446 1336 20480
rect 268 20437 1336 20446
rect 1428 20324 2496 20333
rect 1428 20290 2496 20324
rect 1428 20281 2496 20290
rect 268 20168 1336 20177
rect 268 20134 1336 20168
rect 268 20125 1336 20134
rect 1428 20012 2496 20021
rect 1428 19978 2496 20012
rect 1428 19969 2496 19978
rect 268 19856 1336 19865
rect 268 19822 1336 19856
rect 268 19813 1336 19822
rect 1428 19700 2496 19709
rect 1428 19666 2496 19700
rect 1428 19657 2496 19666
rect 268 19544 1336 19553
rect 268 19510 1336 19544
rect 268 19501 1336 19510
rect 1428 19388 2496 19397
rect 1428 19354 2496 19388
rect 1428 19345 2496 19354
rect 268 19232 1336 19241
rect 268 19198 1336 19232
rect 268 19189 1336 19198
rect 1428 19076 2496 19085
rect 1428 19042 2496 19076
rect 1428 19033 2496 19042
rect 268 18920 1336 18929
rect 268 18886 1336 18920
rect 268 18877 1336 18886
rect 1428 18764 2496 18773
rect 1428 18730 2496 18764
rect 1428 18721 2496 18730
rect 268 18608 1336 18617
rect 268 18574 1336 18608
rect 268 18565 1336 18574
rect 1428 18452 2496 18461
rect 1428 18418 2496 18452
rect 1428 18409 2496 18418
rect 268 18296 1336 18305
rect 268 18262 1336 18296
rect 268 18253 1336 18262
rect 1428 18140 2496 18149
rect 1428 18106 2496 18140
rect 1428 18097 2496 18106
rect 268 17984 1336 17993
rect 268 17950 1336 17984
rect 268 17941 1336 17950
rect 1428 17828 2496 17837
rect 1428 17794 2496 17828
rect 1428 17785 2496 17794
rect 268 17672 1336 17681
rect 268 17638 1336 17672
rect 268 17629 1336 17638
rect 1428 17516 2496 17525
rect 1428 17482 2496 17516
rect 1428 17473 2496 17482
rect 268 17360 1336 17369
rect 268 17326 1336 17360
rect 268 17317 1336 17326
rect 1428 17204 2496 17213
rect 1428 17170 2496 17204
rect 1428 17161 2496 17170
rect 268 17048 1336 17057
rect 268 17014 1336 17048
rect 268 17005 1336 17014
rect 1428 16892 2496 16901
rect 1428 16858 2496 16892
rect 1428 16849 2496 16858
rect 268 16736 1336 16745
rect 268 16702 1336 16736
rect 268 16693 1336 16702
rect 1428 16580 2496 16589
rect 1428 16546 2496 16580
rect 1428 16537 2496 16546
rect 268 16424 1336 16433
rect 268 16390 1336 16424
rect 268 16381 1336 16390
rect 1428 16268 2496 16277
rect 1428 16234 2496 16268
rect 1428 16225 2496 16234
rect 268 16112 1336 16121
rect 268 16078 1336 16112
rect 268 16069 1336 16078
rect 1428 15956 2496 15965
rect 1428 15922 2496 15956
rect 1428 15913 2496 15922
rect 268 15800 1336 15809
rect 268 15766 1336 15800
rect 268 15757 1336 15766
rect 1428 15644 2496 15653
rect 1428 15610 2496 15644
rect 1428 15601 2496 15610
rect 268 15488 1336 15497
rect 268 15454 1336 15488
rect 268 15445 1336 15454
rect 1428 15332 2496 15341
rect 1428 15298 2496 15332
rect 1428 15289 2496 15298
rect 268 15176 1336 15185
rect 268 15142 1336 15176
rect 268 15133 1336 15142
rect 1428 15020 2496 15029
rect 1428 14986 2496 15020
rect 1428 14977 2496 14986
rect 268 14864 1336 14873
rect 268 14830 1336 14864
rect 268 14821 1336 14830
rect 1428 14708 2496 14717
rect 1428 14674 2496 14708
rect 1428 14665 2496 14674
rect 268 14552 1336 14561
rect 268 14518 1336 14552
rect 268 14509 1336 14518
rect 1428 14396 2496 14405
rect 1428 14362 2496 14396
rect 1428 14353 2496 14362
rect 268 14240 1336 14249
rect 268 14206 1336 14240
rect 268 14197 1336 14206
rect 1428 14084 2496 14093
rect 1428 14050 2496 14084
rect 1428 14041 2496 14050
rect 268 13928 1336 13937
rect 268 13894 1336 13928
rect 268 13885 1336 13894
rect 1428 13772 2496 13781
rect 1428 13738 2496 13772
rect 1428 13729 2496 13738
rect 268 13616 1336 13625
rect 268 13582 1336 13616
rect 268 13573 1336 13582
rect 1428 13460 2496 13469
rect 1428 13426 2496 13460
rect 1428 13417 2496 13426
rect 268 13304 1336 13313
rect 268 13270 1336 13304
rect 268 13261 1336 13270
rect 1428 13148 2496 13157
rect 1428 13114 2496 13148
rect 1428 13105 2496 13114
rect 268 12992 1336 13001
rect 268 12958 1336 12992
rect 268 12949 1336 12958
rect 1428 12836 2496 12845
rect 1428 12802 2496 12836
rect 1428 12793 2496 12802
rect 268 12680 1336 12689
rect 268 12646 1336 12680
rect 268 12637 1336 12646
rect 1428 12524 2496 12533
rect 1428 12490 2496 12524
rect 1428 12481 2496 12490
rect 268 12368 1336 12377
rect 268 12334 1336 12368
rect 268 12325 1336 12334
rect 1428 12212 2496 12221
rect 1428 12178 2496 12212
rect 1428 12169 2496 12178
rect 268 12056 1336 12065
rect 268 12022 1336 12056
rect 268 12013 1336 12022
rect 1428 11900 2496 11909
rect 1428 11866 2496 11900
rect 1428 11857 2496 11866
rect 268 11744 1336 11753
rect 268 11710 1336 11744
rect 268 11701 1336 11710
rect 1428 11588 2496 11597
rect 1428 11554 2496 11588
rect 1428 11545 2496 11554
rect 268 11432 1336 11441
rect 268 11398 1336 11432
rect 268 11389 1336 11398
rect 1428 11276 2496 11285
rect 1428 11242 2496 11276
rect 1428 11233 2496 11242
rect 268 11120 1336 11129
rect 268 11086 1336 11120
rect 268 11077 1336 11086
rect 1428 10964 2496 10973
rect 1428 10930 2496 10964
rect 1428 10921 2496 10930
rect 268 10808 1336 10817
rect 268 10774 1336 10808
rect 268 10765 1336 10774
rect 1428 10652 2496 10661
rect 1428 10618 2496 10652
rect 1428 10609 2496 10618
rect 268 10496 1336 10505
rect 268 10462 1336 10496
rect 268 10453 1336 10462
rect 1428 10340 2496 10349
rect 1428 10306 2496 10340
rect 1428 10297 2496 10306
rect 268 10184 1336 10193
rect 268 10150 1336 10184
rect 268 10141 1336 10150
rect 1428 10028 2496 10037
rect 1428 9994 2496 10028
rect 1428 9985 2496 9994
rect 268 9872 1336 9881
rect 268 9838 1336 9872
rect 268 9829 1336 9838
rect 1428 9716 2496 9725
rect 1428 9682 2496 9716
rect 1428 9673 2496 9682
rect 268 9560 1336 9569
rect 268 9526 1336 9560
rect 268 9517 1336 9526
rect 1428 9404 2496 9413
rect 1428 9370 2496 9404
rect 1428 9361 2496 9370
rect 268 9248 1336 9257
rect 268 9214 1336 9248
rect 268 9205 1336 9214
rect 1428 9092 2496 9101
rect 1428 9058 2496 9092
rect 1428 9049 2496 9058
rect 268 8936 1336 8945
rect 268 8902 1336 8936
rect 268 8893 1336 8902
rect 1428 8780 2496 8789
rect 1428 8746 2496 8780
rect 1428 8737 2496 8746
rect 268 8624 1336 8633
rect 268 8590 1336 8624
rect 268 8581 1336 8590
rect 1428 8468 2496 8477
rect 1428 8434 2496 8468
rect 1428 8425 2496 8434
rect 268 8312 1336 8321
rect 268 8278 1336 8312
rect 268 8269 1336 8278
rect 1428 8156 2496 8165
rect 1428 8122 2496 8156
rect 1428 8113 2496 8122
rect 268 8000 1336 8009
rect 268 7966 1336 8000
rect 268 7957 1336 7966
rect 1428 7844 2496 7853
rect 1428 7810 2496 7844
rect 1428 7801 2496 7810
rect 268 7688 1336 7697
rect 268 7654 1336 7688
rect 268 7645 1336 7654
rect 1428 7532 2496 7541
rect 1428 7498 2496 7532
rect 1428 7489 2496 7498
rect 268 7376 1336 7385
rect 268 7342 1336 7376
rect 268 7333 1336 7342
rect 1428 7220 2496 7229
rect 1428 7186 2496 7220
rect 1428 7177 2496 7186
rect 268 7064 1336 7073
rect 268 7030 1336 7064
rect 268 7021 1336 7030
rect 1428 6908 2496 6917
rect 1428 6874 2496 6908
rect 1428 6865 2496 6874
rect 268 6752 1336 6761
rect 268 6718 1336 6752
rect 268 6709 1336 6718
rect 1428 6596 2496 6605
rect 1428 6562 2496 6596
rect 1428 6553 2496 6562
rect 268 6440 1336 6449
rect 268 6406 1336 6440
rect 268 6397 1336 6406
rect 1428 6284 2496 6293
rect 1428 6250 2496 6284
rect 1428 6241 2496 6250
rect 268 6128 1336 6137
rect 268 6094 1336 6128
rect 268 6085 1336 6094
rect 1428 5972 2496 5981
rect 1428 5938 2496 5972
rect 1428 5929 2496 5938
rect 268 5816 1336 5825
rect 268 5782 1336 5816
rect 268 5773 1336 5782
rect 1428 5660 2496 5669
rect 1428 5626 2496 5660
rect 1428 5617 2496 5626
rect 268 5504 1336 5513
rect 268 5470 1336 5504
rect 268 5461 1336 5470
rect 1428 5348 2496 5357
rect 1428 5314 2496 5348
rect 1428 5305 2496 5314
rect 268 5192 1336 5201
rect 268 5158 1336 5192
rect 268 5149 1336 5158
rect 1428 5036 2496 5045
rect 1428 5002 2496 5036
rect 1428 4993 2496 5002
rect 268 4880 1336 4889
rect 268 4846 1336 4880
rect 268 4837 1336 4846
rect 1428 4724 2496 4733
rect 1428 4690 2496 4724
rect 1428 4681 2496 4690
rect 268 4568 1336 4577
rect 268 4534 1336 4568
rect 268 4525 1336 4534
rect 1428 4412 2496 4421
rect 1428 4378 2496 4412
rect 1428 4369 2496 4378
rect 268 4256 1336 4265
rect 268 4222 1336 4256
rect 268 4213 1336 4222
rect 1428 4100 2496 4109
rect 1428 4066 2496 4100
rect 1428 4057 2496 4066
rect 268 3944 1336 3953
rect 268 3910 1336 3944
rect 268 3901 1336 3910
rect 1428 3788 2496 3797
rect 1428 3754 2496 3788
rect 1428 3745 2496 3754
rect 268 3632 1336 3641
rect 268 3598 1336 3632
rect 268 3589 1336 3598
rect 1428 3476 2496 3485
rect 1428 3442 2496 3476
rect 1428 3433 2496 3442
rect 268 3320 1336 3329
rect 268 3286 1336 3320
rect 268 3277 1336 3286
rect 1428 3164 2496 3173
rect 1428 3130 2496 3164
rect 1428 3121 2496 3130
rect 268 3008 1336 3017
rect 268 2974 1336 3008
rect 268 2965 1336 2974
rect 1428 2852 2496 2861
rect 1428 2818 2496 2852
rect 1428 2809 2496 2818
rect 268 2696 1336 2705
rect 268 2662 1336 2696
rect 268 2653 1336 2662
rect 1428 2540 2496 2549
rect 1428 2506 2496 2540
rect 1428 2497 2496 2506
rect 268 2384 1336 2393
rect 268 2350 1336 2384
rect 268 2341 1336 2350
rect 1428 2228 2496 2237
rect 1428 2194 2496 2228
rect 1428 2185 2496 2194
rect 268 2072 1336 2081
rect 268 2038 1336 2072
rect 268 2029 1336 2038
rect 1428 1916 2496 1925
rect 1428 1882 2496 1916
rect 1428 1873 2496 1882
rect 268 1760 1336 1769
rect 268 1726 1336 1760
rect 268 1717 1336 1726
rect 1428 1604 2496 1613
rect 1428 1570 2496 1604
rect 1428 1561 2496 1570
rect 268 1448 1336 1457
rect 268 1414 1336 1448
rect 268 1405 1336 1414
rect 1428 1292 2496 1301
rect 1428 1258 2496 1292
rect 1428 1249 2496 1258
rect 268 1136 1336 1145
rect 268 1102 1336 1136
rect 268 1093 1336 1102
rect 1428 980 2496 989
rect 1428 946 2496 980
rect 1428 937 2496 946
rect 268 824 1336 833
rect 268 790 1336 824
rect 268 781 1336 790
rect 1428 668 2496 677
rect 1428 634 2496 668
rect 1428 625 2496 634
rect 268 512 1336 521
rect 268 478 1336 512
rect 268 469 1336 478
rect 1428 356 2496 365
rect 1428 322 2496 356
rect 1428 313 2496 322
rect 140 233 194 239
rect 268 200 1336 209
rect 268 166 1336 200
rect 268 157 1336 166
<< metal2 >>
rect 262 42901 268 42953
rect 1336 42901 1342 42953
rect 140 42877 194 42883
rect 140 227 194 233
rect 262 42641 1342 42901
rect 262 42589 268 42641
rect 1336 42589 1342 42641
rect 262 42329 1342 42589
rect 262 42277 268 42329
rect 1336 42277 1342 42329
rect 262 42017 1342 42277
rect 262 41965 268 42017
rect 1336 41965 1342 42017
rect 262 41705 1342 41965
rect 262 41653 268 41705
rect 1336 41653 1342 41705
rect 262 41393 1342 41653
rect 262 41341 268 41393
rect 1336 41341 1342 41393
rect 262 41081 1342 41341
rect 262 41029 268 41081
rect 1336 41029 1342 41081
rect 262 40769 1342 41029
rect 262 40717 268 40769
rect 1336 40717 1342 40769
rect 262 40457 1342 40717
rect 262 40405 268 40457
rect 1336 40405 1342 40457
rect 262 40145 1342 40405
rect 262 40093 268 40145
rect 1336 40093 1342 40145
rect 262 39833 1342 40093
rect 262 39781 268 39833
rect 1336 39781 1342 39833
rect 262 39521 1342 39781
rect 262 39469 268 39521
rect 1336 39469 1342 39521
rect 262 39209 1342 39469
rect 262 39157 268 39209
rect 1336 39157 1342 39209
rect 262 38897 1342 39157
rect 262 38845 268 38897
rect 1336 38845 1342 38897
rect 262 38585 1342 38845
rect 262 38533 268 38585
rect 1336 38533 1342 38585
rect 262 38273 1342 38533
rect 262 38221 268 38273
rect 1336 38221 1342 38273
rect 262 37961 1342 38221
rect 262 37909 268 37961
rect 1336 37909 1342 37961
rect 262 37649 1342 37909
rect 262 37597 268 37649
rect 1336 37597 1342 37649
rect 262 37337 1342 37597
rect 262 37285 268 37337
rect 1336 37285 1342 37337
rect 262 37025 1342 37285
rect 262 36973 268 37025
rect 1336 36973 1342 37025
rect 262 36713 1342 36973
rect 262 36661 268 36713
rect 1336 36661 1342 36713
rect 262 36401 1342 36661
rect 262 36349 268 36401
rect 1336 36349 1342 36401
rect 262 36089 1342 36349
rect 262 36037 268 36089
rect 1336 36037 1342 36089
rect 262 35777 1342 36037
rect 262 35725 268 35777
rect 1336 35725 1342 35777
rect 262 35465 1342 35725
rect 262 35413 268 35465
rect 1336 35413 1342 35465
rect 262 35153 1342 35413
rect 262 35101 268 35153
rect 1336 35101 1342 35153
rect 262 34841 1342 35101
rect 262 34789 268 34841
rect 1336 34789 1342 34841
rect 262 34529 1342 34789
rect 262 34477 268 34529
rect 1336 34477 1342 34529
rect 262 34217 1342 34477
rect 262 34165 268 34217
rect 1336 34165 1342 34217
rect 262 33905 1342 34165
rect 262 33853 268 33905
rect 1336 33853 1342 33905
rect 262 33593 1342 33853
rect 262 33541 268 33593
rect 1336 33541 1342 33593
rect 262 33281 1342 33541
rect 262 33229 268 33281
rect 1336 33229 1342 33281
rect 262 32969 1342 33229
rect 262 32917 268 32969
rect 1336 32917 1342 32969
rect 262 32657 1342 32917
rect 262 32605 268 32657
rect 1336 32605 1342 32657
rect 262 32345 1342 32605
rect 262 32293 268 32345
rect 1336 32293 1342 32345
rect 262 32033 1342 32293
rect 262 31981 268 32033
rect 1336 31981 1342 32033
rect 262 31721 1342 31981
rect 262 31669 268 31721
rect 1336 31669 1342 31721
rect 262 31409 1342 31669
rect 262 31357 268 31409
rect 1336 31357 1342 31409
rect 262 31097 1342 31357
rect 262 31045 268 31097
rect 1336 31045 1342 31097
rect 262 30785 1342 31045
rect 262 30733 268 30785
rect 1336 30733 1342 30785
rect 262 30473 1342 30733
rect 262 30421 268 30473
rect 1336 30421 1342 30473
rect 262 30161 1342 30421
rect 262 30109 268 30161
rect 1336 30109 1342 30161
rect 262 29849 1342 30109
rect 262 29797 268 29849
rect 1336 29797 1342 29849
rect 262 29537 1342 29797
rect 262 29485 268 29537
rect 1336 29485 1342 29537
rect 262 29225 1342 29485
rect 262 29173 268 29225
rect 1336 29173 1342 29225
rect 262 28913 1342 29173
rect 262 28861 268 28913
rect 1336 28861 1342 28913
rect 262 28601 1342 28861
rect 262 28549 268 28601
rect 1336 28549 1342 28601
rect 262 28289 1342 28549
rect 262 28237 268 28289
rect 1336 28237 1342 28289
rect 262 27977 1342 28237
rect 262 27925 268 27977
rect 1336 27925 1342 27977
rect 262 27665 1342 27925
rect 262 27613 268 27665
rect 1336 27613 1342 27665
rect 262 27353 1342 27613
rect 262 27301 268 27353
rect 1336 27301 1342 27353
rect 262 27041 1342 27301
rect 262 26989 268 27041
rect 1336 26989 1342 27041
rect 262 26729 1342 26989
rect 262 26677 268 26729
rect 1336 26677 1342 26729
rect 262 26417 1342 26677
rect 262 26365 268 26417
rect 1336 26365 1342 26417
rect 262 26105 1342 26365
rect 262 26053 268 26105
rect 1336 26053 1342 26105
rect 262 25793 1342 26053
rect 262 25741 268 25793
rect 1336 25741 1342 25793
rect 262 25481 1342 25741
rect 262 25429 268 25481
rect 1336 25429 1342 25481
rect 262 25169 1342 25429
rect 262 25117 268 25169
rect 1336 25117 1342 25169
rect 262 24857 1342 25117
rect 262 24805 268 24857
rect 1336 24805 1342 24857
rect 262 24545 1342 24805
rect 262 24493 268 24545
rect 1336 24493 1342 24545
rect 262 24233 1342 24493
rect 262 24181 268 24233
rect 1336 24181 1342 24233
rect 262 23921 1342 24181
rect 262 23869 268 23921
rect 1336 23869 1342 23921
rect 262 23609 1342 23869
rect 262 23557 268 23609
rect 1336 23557 1342 23609
rect 262 23297 1342 23557
rect 262 23245 268 23297
rect 1336 23245 1342 23297
rect 262 22985 1342 23245
rect 262 22933 268 22985
rect 1336 22933 1342 22985
rect 262 22673 1342 22933
rect 262 22621 268 22673
rect 1336 22621 1342 22673
rect 262 22361 1342 22621
rect 262 22309 268 22361
rect 1336 22309 1342 22361
rect 262 22049 1342 22309
rect 262 21997 268 22049
rect 1336 21997 1342 22049
rect 262 21737 1342 21997
rect 262 21685 268 21737
rect 1336 21685 1342 21737
rect 262 21425 1342 21685
rect 262 21373 268 21425
rect 1336 21373 1342 21425
rect 262 21113 1342 21373
rect 262 21061 268 21113
rect 1336 21061 1342 21113
rect 262 20801 1342 21061
rect 262 20749 268 20801
rect 1336 20749 1342 20801
rect 262 20489 1342 20749
rect 262 20437 268 20489
rect 1336 20437 1342 20489
rect 262 20177 1342 20437
rect 262 20125 268 20177
rect 1336 20125 1342 20177
rect 262 19865 1342 20125
rect 262 19813 268 19865
rect 1336 19813 1342 19865
rect 262 19553 1342 19813
rect 262 19501 268 19553
rect 1336 19501 1342 19553
rect 262 19241 1342 19501
rect 262 19189 268 19241
rect 1336 19189 1342 19241
rect 262 18929 1342 19189
rect 262 18877 268 18929
rect 1336 18877 1342 18929
rect 262 18617 1342 18877
rect 262 18565 268 18617
rect 1336 18565 1342 18617
rect 262 18305 1342 18565
rect 262 18253 268 18305
rect 1336 18253 1342 18305
rect 262 17993 1342 18253
rect 262 17941 268 17993
rect 1336 17941 1342 17993
rect 262 17681 1342 17941
rect 262 17629 268 17681
rect 1336 17629 1342 17681
rect 262 17369 1342 17629
rect 262 17317 268 17369
rect 1336 17317 1342 17369
rect 262 17057 1342 17317
rect 262 17005 268 17057
rect 1336 17005 1342 17057
rect 262 16745 1342 17005
rect 262 16693 268 16745
rect 1336 16693 1342 16745
rect 262 16433 1342 16693
rect 262 16381 268 16433
rect 1336 16381 1342 16433
rect 262 16121 1342 16381
rect 262 16069 268 16121
rect 1336 16069 1342 16121
rect 262 15809 1342 16069
rect 262 15757 268 15809
rect 1336 15757 1342 15809
rect 262 15497 1342 15757
rect 262 15445 268 15497
rect 1336 15445 1342 15497
rect 262 15185 1342 15445
rect 262 15133 268 15185
rect 1336 15133 1342 15185
rect 262 14873 1342 15133
rect 262 14821 268 14873
rect 1336 14821 1342 14873
rect 262 14561 1342 14821
rect 262 14509 268 14561
rect 1336 14509 1342 14561
rect 262 14249 1342 14509
rect 262 14197 268 14249
rect 1336 14197 1342 14249
rect 262 13937 1342 14197
rect 262 13885 268 13937
rect 1336 13885 1342 13937
rect 262 13625 1342 13885
rect 262 13573 268 13625
rect 1336 13573 1342 13625
rect 262 13313 1342 13573
rect 262 13261 268 13313
rect 1336 13261 1342 13313
rect 262 13001 1342 13261
rect 262 12949 268 13001
rect 1336 12949 1342 13001
rect 262 12689 1342 12949
rect 262 12637 268 12689
rect 1336 12637 1342 12689
rect 262 12377 1342 12637
rect 262 12325 268 12377
rect 1336 12325 1342 12377
rect 262 12065 1342 12325
rect 262 12013 268 12065
rect 1336 12013 1342 12065
rect 262 11753 1342 12013
rect 262 11701 268 11753
rect 1336 11701 1342 11753
rect 262 11441 1342 11701
rect 262 11389 268 11441
rect 1336 11389 1342 11441
rect 262 11129 1342 11389
rect 262 11077 268 11129
rect 1336 11077 1342 11129
rect 262 10817 1342 11077
rect 262 10765 268 10817
rect 1336 10765 1342 10817
rect 262 10505 1342 10765
rect 262 10453 268 10505
rect 1336 10453 1342 10505
rect 262 10193 1342 10453
rect 262 10141 268 10193
rect 1336 10141 1342 10193
rect 262 9881 1342 10141
rect 262 9829 268 9881
rect 1336 9829 1342 9881
rect 262 9569 1342 9829
rect 262 9517 268 9569
rect 1336 9517 1342 9569
rect 262 9257 1342 9517
rect 262 9205 268 9257
rect 1336 9205 1342 9257
rect 262 8945 1342 9205
rect 262 8893 268 8945
rect 1336 8893 1342 8945
rect 262 8633 1342 8893
rect 262 8581 268 8633
rect 1336 8581 1342 8633
rect 262 8321 1342 8581
rect 262 8269 268 8321
rect 1336 8269 1342 8321
rect 262 8009 1342 8269
rect 262 7957 268 8009
rect 1336 7957 1342 8009
rect 262 7697 1342 7957
rect 262 7645 268 7697
rect 1336 7645 1342 7697
rect 262 7385 1342 7645
rect 262 7333 268 7385
rect 1336 7333 1342 7385
rect 262 7073 1342 7333
rect 262 7021 268 7073
rect 1336 7021 1342 7073
rect 262 6761 1342 7021
rect 262 6709 268 6761
rect 1336 6709 1342 6761
rect 262 6449 1342 6709
rect 262 6397 268 6449
rect 1336 6397 1342 6449
rect 262 6137 1342 6397
rect 262 6085 268 6137
rect 1336 6085 1342 6137
rect 262 5825 1342 6085
rect 262 5773 268 5825
rect 1336 5773 1342 5825
rect 262 5513 1342 5773
rect 262 5461 268 5513
rect 1336 5461 1342 5513
rect 262 5201 1342 5461
rect 262 5149 268 5201
rect 1336 5149 1342 5201
rect 262 4889 1342 5149
rect 262 4837 268 4889
rect 1336 4837 1342 4889
rect 262 4577 1342 4837
rect 262 4525 268 4577
rect 1336 4525 1342 4577
rect 262 4265 1342 4525
rect 262 4213 268 4265
rect 1336 4213 1342 4265
rect 262 3953 1342 4213
rect 262 3901 268 3953
rect 1336 3901 1342 3953
rect 262 3641 1342 3901
rect 262 3589 268 3641
rect 1336 3589 1342 3641
rect 262 3329 1342 3589
rect 262 3277 268 3329
rect 1336 3277 1342 3329
rect 262 3017 1342 3277
rect 262 2965 268 3017
rect 1336 2965 1342 3017
rect 262 2705 1342 2965
rect 262 2653 268 2705
rect 1336 2653 1342 2705
rect 262 2393 1342 2653
rect 262 2341 268 2393
rect 1336 2341 1342 2393
rect 262 2081 1342 2341
rect 262 2029 268 2081
rect 1336 2029 1342 2081
rect 262 1769 1342 2029
rect 262 1717 268 1769
rect 1336 1717 1342 1769
rect 262 1457 1342 1717
rect 262 1405 268 1457
rect 1336 1405 1342 1457
rect 262 1145 1342 1405
rect 262 1093 268 1145
rect 1336 1093 1342 1145
rect 262 833 1342 1093
rect 262 781 268 833
rect 1336 781 1342 833
rect 262 521 1342 781
rect 262 469 268 521
rect 1336 469 1342 521
rect 262 209 1342 469
rect 262 157 268 209
rect 1336 157 1342 209
rect 1422 42797 2502 42953
rect 1422 42745 1428 42797
rect 2496 42745 2502 42797
rect 1422 42485 2502 42745
rect 1422 42433 1428 42485
rect 2496 42433 2502 42485
rect 1422 42173 2502 42433
rect 1422 42121 1428 42173
rect 2496 42121 2502 42173
rect 1422 41861 2502 42121
rect 1422 41809 1428 41861
rect 2496 41809 2502 41861
rect 1422 41549 2502 41809
rect 1422 41497 1428 41549
rect 2496 41497 2502 41549
rect 1422 41237 2502 41497
rect 1422 41185 1428 41237
rect 2496 41185 2502 41237
rect 1422 40925 2502 41185
rect 1422 40873 1428 40925
rect 2496 40873 2502 40925
rect 1422 40613 2502 40873
rect 1422 40561 1428 40613
rect 2496 40561 2502 40613
rect 1422 40301 2502 40561
rect 1422 40249 1428 40301
rect 2496 40249 2502 40301
rect 1422 39989 2502 40249
rect 1422 39937 1428 39989
rect 2496 39937 2502 39989
rect 1422 39677 2502 39937
rect 1422 39625 1428 39677
rect 2496 39625 2502 39677
rect 1422 39365 2502 39625
rect 1422 39313 1428 39365
rect 2496 39313 2502 39365
rect 1422 39053 2502 39313
rect 1422 39001 1428 39053
rect 2496 39001 2502 39053
rect 1422 38741 2502 39001
rect 1422 38689 1428 38741
rect 2496 38689 2502 38741
rect 1422 38429 2502 38689
rect 1422 38377 1428 38429
rect 2496 38377 2502 38429
rect 1422 38117 2502 38377
rect 1422 38065 1428 38117
rect 2496 38065 2502 38117
rect 1422 37805 2502 38065
rect 1422 37753 1428 37805
rect 2496 37753 2502 37805
rect 1422 37493 2502 37753
rect 1422 37441 1428 37493
rect 2496 37441 2502 37493
rect 1422 37181 2502 37441
rect 1422 37129 1428 37181
rect 2496 37129 2502 37181
rect 1422 36869 2502 37129
rect 1422 36817 1428 36869
rect 2496 36817 2502 36869
rect 1422 36557 2502 36817
rect 1422 36505 1428 36557
rect 2496 36505 2502 36557
rect 1422 36245 2502 36505
rect 1422 36193 1428 36245
rect 2496 36193 2502 36245
rect 1422 35933 2502 36193
rect 1422 35881 1428 35933
rect 2496 35881 2502 35933
rect 1422 35621 2502 35881
rect 1422 35569 1428 35621
rect 2496 35569 2502 35621
rect 1422 35309 2502 35569
rect 1422 35257 1428 35309
rect 2496 35257 2502 35309
rect 1422 34997 2502 35257
rect 1422 34945 1428 34997
rect 2496 34945 2502 34997
rect 1422 34685 2502 34945
rect 1422 34633 1428 34685
rect 2496 34633 2502 34685
rect 1422 34373 2502 34633
rect 1422 34321 1428 34373
rect 2496 34321 2502 34373
rect 1422 34061 2502 34321
rect 1422 34009 1428 34061
rect 2496 34009 2502 34061
rect 1422 33749 2502 34009
rect 1422 33697 1428 33749
rect 2496 33697 2502 33749
rect 1422 33437 2502 33697
rect 1422 33385 1428 33437
rect 2496 33385 2502 33437
rect 1422 33125 2502 33385
rect 1422 33073 1428 33125
rect 2496 33073 2502 33125
rect 1422 32813 2502 33073
rect 1422 32761 1428 32813
rect 2496 32761 2502 32813
rect 1422 32501 2502 32761
rect 1422 32449 1428 32501
rect 2496 32449 2502 32501
rect 1422 32189 2502 32449
rect 1422 32137 1428 32189
rect 2496 32137 2502 32189
rect 1422 31877 2502 32137
rect 1422 31825 1428 31877
rect 2496 31825 2502 31877
rect 1422 31565 2502 31825
rect 1422 31513 1428 31565
rect 2496 31513 2502 31565
rect 1422 31253 2502 31513
rect 1422 31201 1428 31253
rect 2496 31201 2502 31253
rect 1422 30941 2502 31201
rect 1422 30889 1428 30941
rect 2496 30889 2502 30941
rect 1422 30629 2502 30889
rect 1422 30577 1428 30629
rect 2496 30577 2502 30629
rect 1422 30317 2502 30577
rect 1422 30265 1428 30317
rect 2496 30265 2502 30317
rect 1422 30005 2502 30265
rect 1422 29953 1428 30005
rect 2496 29953 2502 30005
rect 1422 29693 2502 29953
rect 1422 29641 1428 29693
rect 2496 29641 2502 29693
rect 1422 29381 2502 29641
rect 1422 29329 1428 29381
rect 2496 29329 2502 29381
rect 1422 29069 2502 29329
rect 1422 29017 1428 29069
rect 2496 29017 2502 29069
rect 1422 28757 2502 29017
rect 1422 28705 1428 28757
rect 2496 28705 2502 28757
rect 1422 28445 2502 28705
rect 1422 28393 1428 28445
rect 2496 28393 2502 28445
rect 1422 28133 2502 28393
rect 1422 28081 1428 28133
rect 2496 28081 2502 28133
rect 1422 27821 2502 28081
rect 1422 27769 1428 27821
rect 2496 27769 2502 27821
rect 1422 27509 2502 27769
rect 1422 27457 1428 27509
rect 2496 27457 2502 27509
rect 1422 27197 2502 27457
rect 1422 27145 1428 27197
rect 2496 27145 2502 27197
rect 1422 26885 2502 27145
rect 1422 26833 1428 26885
rect 2496 26833 2502 26885
rect 1422 26573 2502 26833
rect 1422 26521 1428 26573
rect 2496 26521 2502 26573
rect 1422 26261 2502 26521
rect 1422 26209 1428 26261
rect 2496 26209 2502 26261
rect 1422 25949 2502 26209
rect 1422 25897 1428 25949
rect 2496 25897 2502 25949
rect 1422 25637 2502 25897
rect 1422 25585 1428 25637
rect 2496 25585 2502 25637
rect 1422 25325 2502 25585
rect 1422 25273 1428 25325
rect 2496 25273 2502 25325
rect 1422 25013 2502 25273
rect 1422 24961 1428 25013
rect 2496 24961 2502 25013
rect 1422 24701 2502 24961
rect 1422 24649 1428 24701
rect 2496 24649 2502 24701
rect 1422 24389 2502 24649
rect 1422 24337 1428 24389
rect 2496 24337 2502 24389
rect 1422 24077 2502 24337
rect 1422 24025 1428 24077
rect 2496 24025 2502 24077
rect 1422 23765 2502 24025
rect 1422 23713 1428 23765
rect 2496 23713 2502 23765
rect 1422 23453 2502 23713
rect 1422 23401 1428 23453
rect 2496 23401 2502 23453
rect 1422 23141 2502 23401
rect 1422 23089 1428 23141
rect 2496 23089 2502 23141
rect 1422 22829 2502 23089
rect 1422 22777 1428 22829
rect 2496 22777 2502 22829
rect 1422 22517 2502 22777
rect 1422 22465 1428 22517
rect 2496 22465 2502 22517
rect 1422 22205 2502 22465
rect 1422 22153 1428 22205
rect 2496 22153 2502 22205
rect 1422 21893 2502 22153
rect 1422 21841 1428 21893
rect 2496 21841 2502 21893
rect 1422 21581 2502 21841
rect 1422 21529 1428 21581
rect 2496 21529 2502 21581
rect 1422 21269 2502 21529
rect 1422 21217 1428 21269
rect 2496 21217 2502 21269
rect 1422 20957 2502 21217
rect 1422 20905 1428 20957
rect 2496 20905 2502 20957
rect 1422 20645 2502 20905
rect 1422 20593 1428 20645
rect 2496 20593 2502 20645
rect 1422 20333 2502 20593
rect 1422 20281 1428 20333
rect 2496 20281 2502 20333
rect 1422 20021 2502 20281
rect 1422 19969 1428 20021
rect 2496 19969 2502 20021
rect 1422 19709 2502 19969
rect 1422 19657 1428 19709
rect 2496 19657 2502 19709
rect 1422 19397 2502 19657
rect 1422 19345 1428 19397
rect 2496 19345 2502 19397
rect 1422 19085 2502 19345
rect 1422 19033 1428 19085
rect 2496 19033 2502 19085
rect 1422 18773 2502 19033
rect 1422 18721 1428 18773
rect 2496 18721 2502 18773
rect 1422 18461 2502 18721
rect 1422 18409 1428 18461
rect 2496 18409 2502 18461
rect 1422 18149 2502 18409
rect 1422 18097 1428 18149
rect 2496 18097 2502 18149
rect 1422 17837 2502 18097
rect 1422 17785 1428 17837
rect 2496 17785 2502 17837
rect 1422 17525 2502 17785
rect 1422 17473 1428 17525
rect 2496 17473 2502 17525
rect 1422 17213 2502 17473
rect 1422 17161 1428 17213
rect 2496 17161 2502 17213
rect 1422 16901 2502 17161
rect 1422 16849 1428 16901
rect 2496 16849 2502 16901
rect 1422 16589 2502 16849
rect 1422 16537 1428 16589
rect 2496 16537 2502 16589
rect 1422 16277 2502 16537
rect 1422 16225 1428 16277
rect 2496 16225 2502 16277
rect 1422 15965 2502 16225
rect 1422 15913 1428 15965
rect 2496 15913 2502 15965
rect 1422 15653 2502 15913
rect 1422 15601 1428 15653
rect 2496 15601 2502 15653
rect 1422 15341 2502 15601
rect 1422 15289 1428 15341
rect 2496 15289 2502 15341
rect 1422 15029 2502 15289
rect 1422 14977 1428 15029
rect 2496 14977 2502 15029
rect 1422 14717 2502 14977
rect 1422 14665 1428 14717
rect 2496 14665 2502 14717
rect 1422 14405 2502 14665
rect 1422 14353 1428 14405
rect 2496 14353 2502 14405
rect 1422 14093 2502 14353
rect 1422 14041 1428 14093
rect 2496 14041 2502 14093
rect 1422 13781 2502 14041
rect 1422 13729 1428 13781
rect 2496 13729 2502 13781
rect 1422 13469 2502 13729
rect 1422 13417 1428 13469
rect 2496 13417 2502 13469
rect 1422 13157 2502 13417
rect 1422 13105 1428 13157
rect 2496 13105 2502 13157
rect 1422 12845 2502 13105
rect 1422 12793 1428 12845
rect 2496 12793 2502 12845
rect 1422 12533 2502 12793
rect 1422 12481 1428 12533
rect 2496 12481 2502 12533
rect 1422 12221 2502 12481
rect 1422 12169 1428 12221
rect 2496 12169 2502 12221
rect 1422 11909 2502 12169
rect 1422 11857 1428 11909
rect 2496 11857 2502 11909
rect 1422 11597 2502 11857
rect 1422 11545 1428 11597
rect 2496 11545 2502 11597
rect 1422 11285 2502 11545
rect 1422 11233 1428 11285
rect 2496 11233 2502 11285
rect 1422 10973 2502 11233
rect 1422 10921 1428 10973
rect 2496 10921 2502 10973
rect 1422 10661 2502 10921
rect 1422 10609 1428 10661
rect 2496 10609 2502 10661
rect 1422 10349 2502 10609
rect 1422 10297 1428 10349
rect 2496 10297 2502 10349
rect 1422 10037 2502 10297
rect 1422 9985 1428 10037
rect 2496 9985 2502 10037
rect 1422 9725 2502 9985
rect 1422 9673 1428 9725
rect 2496 9673 2502 9725
rect 1422 9413 2502 9673
rect 1422 9361 1428 9413
rect 2496 9361 2502 9413
rect 1422 9101 2502 9361
rect 1422 9049 1428 9101
rect 2496 9049 2502 9101
rect 1422 8789 2502 9049
rect 1422 8737 1428 8789
rect 2496 8737 2502 8789
rect 1422 8477 2502 8737
rect 1422 8425 1428 8477
rect 2496 8425 2502 8477
rect 1422 8165 2502 8425
rect 1422 8113 1428 8165
rect 2496 8113 2502 8165
rect 1422 7853 2502 8113
rect 1422 7801 1428 7853
rect 2496 7801 2502 7853
rect 1422 7541 2502 7801
rect 1422 7489 1428 7541
rect 2496 7489 2502 7541
rect 1422 7229 2502 7489
rect 1422 7177 1428 7229
rect 2496 7177 2502 7229
rect 1422 6917 2502 7177
rect 1422 6865 1428 6917
rect 2496 6865 2502 6917
rect 1422 6605 2502 6865
rect 1422 6553 1428 6605
rect 2496 6553 2502 6605
rect 1422 6293 2502 6553
rect 1422 6241 1428 6293
rect 2496 6241 2502 6293
rect 1422 5981 2502 6241
rect 1422 5929 1428 5981
rect 2496 5929 2502 5981
rect 1422 5669 2502 5929
rect 1422 5617 1428 5669
rect 2496 5617 2502 5669
rect 1422 5357 2502 5617
rect 1422 5305 1428 5357
rect 2496 5305 2502 5357
rect 1422 5045 2502 5305
rect 1422 4993 1428 5045
rect 2496 4993 2502 5045
rect 1422 4733 2502 4993
rect 1422 4681 1428 4733
rect 2496 4681 2502 4733
rect 1422 4421 2502 4681
rect 1422 4369 1428 4421
rect 2496 4369 2502 4421
rect 1422 4109 2502 4369
rect 1422 4057 1428 4109
rect 2496 4057 2502 4109
rect 1422 3797 2502 4057
rect 1422 3745 1428 3797
rect 2496 3745 2502 3797
rect 1422 3485 2502 3745
rect 1422 3433 1428 3485
rect 2496 3433 2502 3485
rect 1422 3173 2502 3433
rect 1422 3121 1428 3173
rect 2496 3121 2502 3173
rect 1422 2861 2502 3121
rect 1422 2809 1428 2861
rect 2496 2809 2502 2861
rect 1422 2549 2502 2809
rect 1422 2497 1428 2549
rect 2496 2497 2502 2549
rect 1422 2237 2502 2497
rect 1422 2185 1428 2237
rect 2496 2185 2502 2237
rect 1422 1925 2502 2185
rect 1422 1873 1428 1925
rect 2496 1873 2502 1925
rect 1422 1613 2502 1873
rect 1422 1561 1428 1613
rect 2496 1561 2502 1613
rect 1422 1301 2502 1561
rect 1422 1249 1428 1301
rect 2496 1249 2502 1301
rect 1422 989 2502 1249
rect 1422 937 1428 989
rect 2496 937 2502 989
rect 1422 677 2502 937
rect 1422 625 1428 677
rect 2496 625 2502 677
rect 1422 365 2502 625
rect 1422 313 1428 365
rect 2496 313 2502 365
rect 1422 157 2502 313
<< end >>
